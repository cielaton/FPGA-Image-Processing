`include "parameter.v"

module image_read();
endmodule
