//`include "parameter.v"
module image_read #(
parameter WIDTH = 40, HEIGHT = 20,
    STARTUP_DELAY = 100,  //Delay during startup time
    HSYNC_DELAY = 160,  //Hsync pulse delay
    BRIGHTNESS_VALUE = 100,  //For brightness operation
    THRESHOLD = 90,  //For threshold operation
    SIGN = 1  /*
              For brightness operation.
              SIGN = 0 -> Brightness subtraction
              SIGN = 1 -> Brightness addition
              */
) (
    input HCLK,  // Clock
    input HRESET,  // Reset (active low)
    output VSYNC,  // Indicate whether the entire image is transmitted
    output reg HSYNC,  // Indicate whether one line of the image is transmitted

    output reg [7:0] DATA_R0,  // 8 bit Red data (even)
    output reg [7:0] DATA_G0,  // 8 bit Green data (even)
    output reg [7:0] DATA_B0,  // 8 bit Blue data (even)
    output reg [7:0] DATA_R1,  // 8 bit Red data (odd)
    output reg [7:0] DATA_G1,  // 8 bit Green data (odd)
    output reg [7:0] DATA_B1,  // 8 bit Blue data (odd)
    // We will process and transmit 2 pixels in parallel for faster processing
    output ctrl_done,  // Done flag

    input increaseBrightness,
    input decreaseBrightness,
    input threshold,
    input invert,
    output started
);

  parameter sizeOfWidth = 8;  // Data width
  parameter imageDataLenght = WIDTH * HEIGHT * 3;  // Lenght in bytes, each byte represent one of Red, Green, Blue value

  // local parameters for FSM
  localparam ST_IDLE = 2'b00;  // Idle state
  localparam ST_VSYNC = 2'b01;  // State for creating vsync
  localparam ST_HSYNC = 2'b10;  // State for creating hsync
  localparam ST_DATA = 2'b11;  // State for data processing

  reg [1:0] currentState, nextState;
  reg start;  // Signal the FSM begin to operate
  reg HRESETDelay;  // Use to create start signal
  reg vsyncControlSignal, hsyncControlSignal;
  reg [8:0] vsyncControlCounter, hsyncControlCounter;
  reg dataProcessingControlSignal;

  reg [7:0] totalMemory[0:imageDataLenght - 1];  // Memory to store 8-bit data image 

  // Temporary memory to save image data
  integer tempBMP[0:imageDataLenght - 1];
  integer tempRedValue[0:WIDTH * HEIGHT - 1];
  integer tempGreenValue[0:WIDTH * HEIGHT - 1];
  integer tempBlueValue[0:WIDTH * HEIGHT - 1];

  integer i, j;  // Counting variables

  integer
      tempConBriR0,
      tempConBriR1,
      tempConBriG0,
      tempConBriG1,
      tempConBriB0,
      tempConBriB1;  // Temporary variables in contrast and brightness operation

  integer
      tempInvThre,
      tempInvThre1,
      tempInvThre2,
      tempInvThre4;  // Temporary variables in invert and threshold operation

  reg [ 9:0] rowIndex;
  reg [10:0] colIndex;
  reg [18:0] pixelDataCount;  // For creating the done flag

  assign started = start;

  // --- READING IMAGE ---
initial begin
totalMemory[0] = 8'hf2;totalMemory[1] = 8'hcd;totalMemory[2] = 8'hd1;totalMemory[3] = 8'hf4;totalMemory[4] = 8'hd3;totalMemory[5] = 8'hd5;totalMemory[6] = 8'hf7;totalMemory[7] = 8'hd7;totalMemory[8] = 8'hda;totalMemory[9] = 8'hfb;totalMemory[10] = 8'hdd;totalMemory[11] = 8'he0;totalMemory[12] = 8'hfe;totalMemory[13] = 8'he6;totalMemory[14] = 8'he9;totalMemory[15] = 8'hfe;totalMemory[16] = 8'he4;totalMemory[17] = 8'he8;totalMemory[18] = 8'hfa;totalMemory[19] = 8'hdc;totalMemory[20] = 8'hdf;totalMemory[21] = 8'hfa;totalMemory[22] = 8'hd8;totalMemory[23] = 8'hda;totalMemory[24] = 8'hfb;totalMemory[25] = 8'hd9;totalMemory[26] = 8'hda;totalMemory[27] = 8'hfd;totalMemory[28] = 8'hd9;totalMemory[29] = 8'hd8;totalMemory[30] = 8'hff;totalMemory[31] = 8'hda;totalMemory[32] = 8'hd6;totalMemory[33] = 8'hff;totalMemory[34] = 8'he0;totalMemory[35] = 8'hdb;totalMemory[36] = 8'hff;totalMemory[37] = 8'he8;totalMemory[38] = 8'he2;totalMemory[39] = 8'hff;totalMemory[40] = 8'he9;totalMemory[41] = 8'he4;totalMemory[42] = 8'hff;totalMemory[43] = 8'he6;totalMemory[44] = 8'he0;totalMemory[45] = 8'hff;totalMemory[46] = 8'he7;totalMemory[47] = 8'he1;totalMemory[48] = 8'hfa;totalMemory[49] = 8'he6;totalMemory[50] = 8'he0;totalMemory[51] = 8'hc1;totalMemory[52] = 8'hb0;totalMemory[53] = 8'hab;totalMemory[54] = 8'h6b;totalMemory[55] = 8'h5e;totalMemory[56] = 8'h55;totalMemory[57] = 8'h3c;totalMemory[58] = 8'h34;totalMemory[59] = 8'h25;totalMemory[60] = 8'h3b;totalMemory[61] = 8'h36;totalMemory[62] = 8'h18;totalMemory[63] = 8'h55;totalMemory[64] = 8'h50;totalMemory[65] = 8'h1a;totalMemory[66] = 8'h77;totalMemory[67] = 8'h6d;totalMemory[68] = 8'h1f;totalMemory[69] = 8'h96;totalMemory[70] = 8'h83;totalMemory[71] = 8'h1d;totalMemory[72] = 8'hae;totalMemory[73] = 8'h94;totalMemory[74] = 8'h1d;totalMemory[75] = 8'hbb;totalMemory[76] = 8'h9a;totalMemory[77] = 8'h1a;totalMemory[78] = 8'hbc;totalMemory[79] = 8'h98;totalMemory[80] = 8'h13;totalMemory[81] = 8'hba;totalMemory[82] = 8'h96;totalMemory[83] = 8'hf;totalMemory[84] = 8'hbe;totalMemory[85] = 8'h98;totalMemory[86] = 8'hd;totalMemory[87] = 8'hca;totalMemory[88] = 8'h9f;totalMemory[89] = 8'hc;totalMemory[90] = 8'hd3;totalMemory[91] = 8'ha5;totalMemory[92] = 8'hb;totalMemory[93] = 8'hd4;totalMemory[94] = 8'ha5;totalMemory[95] = 8'h6;totalMemory[96] = 8'hd5;totalMemory[97] = 8'ha5;totalMemory[98] = 8'h2;totalMemory[99] = 8'hd7;totalMemory[100] = 8'ha4;totalMemory[101] = 8'h0;totalMemory[102] = 8'hdb;totalMemory[103] = 8'ha7;totalMemory[104] = 8'h0;totalMemory[105] = 8'he2;totalMemory[106] = 8'hae;totalMemory[107] = 8'h0;totalMemory[108] = 8'he5;totalMemory[109] = 8'hb2;totalMemory[110] = 8'h0;totalMemory[111] = 8'he6;totalMemory[112] = 8'hb1;totalMemory[113] = 8'h0;totalMemory[114] = 8'he8;totalMemory[115] = 8'hb2;totalMemory[116] = 8'h0;totalMemory[117] = 8'he9;totalMemory[118] = 8'hb4;totalMemory[119] = 8'h0;totalMemory[120] = 8'hf5;totalMemory[121] = 8'hcf;totalMemory[122] = 8'hd2;totalMemory[123] = 8'hfc;totalMemory[124] = 8'hdd;totalMemory[125] = 8'hde;totalMemory[126] = 8'hff;totalMemory[127] = 8'he6;totalMemory[128] = 8'he7;totalMemory[129] = 8'hfe;totalMemory[130] = 8'he5;totalMemory[131] = 8'he9;totalMemory[132] = 8'hfe;totalMemory[133] = 8'he5;totalMemory[134] = 8'hea;totalMemory[135] = 8'hff;totalMemory[136] = 8'he7;totalMemory[137] = 8'hec;totalMemory[138] = 8'hff;totalMemory[139] = 8'he6;totalMemory[140] = 8'he9;totalMemory[141] = 8'hff;totalMemory[142] = 8'he4;totalMemory[143] = 8'he6;totalMemory[144] = 8'hff;totalMemory[145] = 8'he5;totalMemory[146] = 8'he4;totalMemory[147] = 8'hff;totalMemory[148] = 8'he4;totalMemory[149] = 8'he2;totalMemory[150] = 8'hff;totalMemory[151] = 8'he3;totalMemory[152] = 8'hde;totalMemory[153] = 8'hff;totalMemory[154] = 8'he4;totalMemory[155] = 8'hdf;totalMemory[156] = 8'hff;totalMemory[157] = 8'he6;totalMemory[158] = 8'he1;totalMemory[159] = 8'hff;totalMemory[160] = 8'hec;totalMemory[161] = 8'he5;totalMemory[162] = 8'hff;totalMemory[163] = 8'hed;totalMemory[164] = 8'he6;totalMemory[165] = 8'hff;totalMemory[166] = 8'hee;totalMemory[167] = 8'he8;totalMemory[168] = 8'he3;totalMemory[169] = 8'hd3;totalMemory[170] = 8'hcc;totalMemory[171] = 8'h92;totalMemory[172] = 8'h84;totalMemory[173] = 8'h7d;totalMemory[174] = 8'h4a;totalMemory[175] = 8'h40;totalMemory[176] = 8'h33;totalMemory[177] = 8'h35;totalMemory[178] = 8'h2e;totalMemory[179] = 8'h18;totalMemory[180] = 8'h4a;totalMemory[181] = 8'h42;totalMemory[182] = 8'h19;totalMemory[183] = 8'h70;totalMemory[184] = 8'h66;totalMemory[185] = 8'h20;totalMemory[186] = 8'h91;totalMemory[187] = 8'h80;totalMemory[188] = 8'h22;totalMemory[189] = 8'ha7;totalMemory[190] = 8'h8e;totalMemory[191] = 8'h1d;totalMemory[192] = 8'hb4;totalMemory[193] = 8'h96;totalMemory[194] = 8'h1b;totalMemory[195] = 8'hb6;totalMemory[196] = 8'h96;totalMemory[197] = 8'h18;totalMemory[198] = 8'hb0;totalMemory[199] = 8'h8f;totalMemory[200] = 8'h10;totalMemory[201] = 8'hb0;totalMemory[202] = 8'h8e;totalMemory[203] = 8'hd;totalMemory[204] = 8'hbc;totalMemory[205] = 8'h98;totalMemory[206] = 8'h10;totalMemory[207] = 8'hc9;totalMemory[208] = 8'h9f;totalMemory[209] = 8'he;totalMemory[210] = 8'hcf;totalMemory[211] = 8'ha2;totalMemory[212] = 8'h9;totalMemory[213] = 8'hd0;totalMemory[214] = 8'ha2;totalMemory[215] = 8'h4;totalMemory[216] = 8'hd2;totalMemory[217] = 8'ha3;totalMemory[218] = 8'h1;totalMemory[219] = 8'hd8;totalMemory[220] = 8'ha8;totalMemory[221] = 8'h2;totalMemory[222] = 8'he0;totalMemory[223] = 8'hae;totalMemory[224] = 8'h2;totalMemory[225] = 8'he5;totalMemory[226] = 8'hb2;totalMemory[227] = 8'h1;totalMemory[228] = 8'he7;totalMemory[229] = 8'hb3;totalMemory[230] = 8'h0;totalMemory[231] = 8'he8;totalMemory[232] = 8'hb4;totalMemory[233] = 8'h0;totalMemory[234] = 8'he9;totalMemory[235] = 8'hb5;totalMemory[236] = 8'h0;totalMemory[237] = 8'he7;totalMemory[238] = 8'hb4;totalMemory[239] = 8'h0;totalMemory[240] = 8'hf1;totalMemory[241] = 8'hca;totalMemory[242] = 8'hce;totalMemory[243] = 8'hf3;totalMemory[244] = 8'hd0;totalMemory[245] = 8'hd2;totalMemory[246] = 8'hf8;totalMemory[247] = 8'hdb;totalMemory[248] = 8'hdc;totalMemory[249] = 8'hfd;totalMemory[250] = 8'he2;totalMemory[251] = 8'he5;totalMemory[252] = 8'hff;totalMemory[253] = 8'he2;totalMemory[254] = 8'he6;totalMemory[255] = 8'hff;totalMemory[256] = 8'he4;totalMemory[257] = 8'he8;totalMemory[258] = 8'hff;totalMemory[259] = 8'he5;totalMemory[260] = 8'he8;totalMemory[261] = 8'hff;totalMemory[262] = 8'he3;totalMemory[263] = 8'he3;totalMemory[264] = 8'hff;totalMemory[265] = 8'he1;totalMemory[266] = 8'he0;totalMemory[267] = 8'hff;totalMemory[268] = 8'he5;totalMemory[269] = 8'he1;totalMemory[270] = 8'hff;totalMemory[271] = 8'he7;totalMemory[272] = 8'he2;totalMemory[273] = 8'hff;totalMemory[274] = 8'he6;totalMemory[275] = 8'he1;totalMemory[276] = 8'hff;totalMemory[277] = 8'he4;totalMemory[278] = 8'hdf;totalMemory[279] = 8'hff;totalMemory[280] = 8'hea;totalMemory[281] = 8'he5;totalMemory[282] = 8'hff;totalMemory[283] = 8'hf2;totalMemory[284] = 8'hed;totalMemory[285] = 8'hf1;totalMemory[286] = 8'he4;totalMemory[287] = 8'he0;totalMemory[288] = 8'hb0;totalMemory[289] = 8'ha3;totalMemory[290] = 8'h9e;totalMemory[291] = 8'h5f;totalMemory[292] = 8'h56;totalMemory[293] = 8'h4c;totalMemory[294] = 8'h38;totalMemory[295] = 8'h31;totalMemory[296] = 8'h1d;totalMemory[297] = 8'h3f;totalMemory[298] = 8'h38;totalMemory[299] = 8'h14;totalMemory[300] = 8'h65;totalMemory[301] = 8'h5a;totalMemory[302] = 8'h1e;totalMemory[303] = 8'h8e;totalMemory[304] = 8'h7c;totalMemory[305] = 8'h23;totalMemory[306] = 8'ha9;totalMemory[307] = 8'h8f;totalMemory[308] = 8'h22;totalMemory[309] = 8'hb4;totalMemory[310] = 8'h96;totalMemory[311] = 8'h1e;totalMemory[312] = 8'hb1;totalMemory[313] = 8'h93;totalMemory[314] = 8'h1a;totalMemory[315] = 8'ha4;totalMemory[316] = 8'h8b;totalMemory[317] = 8'h16;totalMemory[318] = 8'h9f;totalMemory[319] = 8'h85;totalMemory[320] = 8'hf;totalMemory[321] = 8'had;totalMemory[322] = 8'h8d;totalMemory[323] = 8'hf;totalMemory[324] = 8'hc0;totalMemory[325] = 8'h9c;totalMemory[326] = 8'h13;totalMemory[327] = 8'hc9;totalMemory[328] = 8'ha0;totalMemory[329] = 8'h10;totalMemory[330] = 8'hca;totalMemory[331] = 8'h9e;totalMemory[332] = 8'h8;totalMemory[333] = 8'hcc;totalMemory[334] = 8'h9e;totalMemory[335] = 8'h7;totalMemory[336] = 8'hd3;totalMemory[337] = 8'ha4;totalMemory[338] = 8'h7;totalMemory[339] = 8'hdd;totalMemory[340] = 8'had;totalMemory[341] = 8'h8;totalMemory[342] = 8'he4;totalMemory[343] = 8'hb2;totalMemory[344] = 8'h5;totalMemory[345] = 8'he6;totalMemory[346] = 8'hb2;totalMemory[347] = 8'h1;totalMemory[348] = 8'he6;totalMemory[349] = 8'hb2;totalMemory[350] = 8'h0;totalMemory[351] = 8'he7;totalMemory[352] = 8'hb3;totalMemory[353] = 8'h0;totalMemory[354] = 8'he6;totalMemory[355] = 8'hb3;totalMemory[356] = 8'h0;totalMemory[357] = 8'he3;totalMemory[358] = 8'hb1;totalMemory[359] = 8'h0;totalMemory[360] = 8'hec;totalMemory[361] = 8'hc7;totalMemory[362] = 8'hca;totalMemory[363] = 8'hee;totalMemory[364] = 8'hc6;totalMemory[365] = 8'hc9;totalMemory[366] = 8'hf1;totalMemory[367] = 8'hc9;totalMemory[368] = 8'hcb;totalMemory[369] = 8'hf7;totalMemory[370] = 8'hd1;totalMemory[371] = 8'hd3;totalMemory[372] = 8'hfc;totalMemory[373] = 8'hd9;totalMemory[374] = 8'hdb;totalMemory[375] = 8'hff;totalMemory[376] = 8'he1;totalMemory[377] = 8'he4;totalMemory[378] = 8'hff;totalMemory[379] = 8'he6;totalMemory[380] = 8'he8;totalMemory[381] = 8'hff;totalMemory[382] = 8'he3;totalMemory[383] = 8'he4;totalMemory[384] = 8'hff;totalMemory[385] = 8'he0;totalMemory[386] = 8'hde;totalMemory[387] = 8'hff;totalMemory[388] = 8'he3;totalMemory[389] = 8'hde;totalMemory[390] = 8'hff;totalMemory[391] = 8'he7;totalMemory[392] = 8'he2;totalMemory[393] = 8'hff;totalMemory[394] = 8'heb;totalMemory[395] = 8'he6;totalMemory[396] = 8'hff;totalMemory[397] = 8'hee;totalMemory[398] = 8'hea;totalMemory[399] = 8'hff;totalMemory[400] = 8'hf5;totalMemory[401] = 8'hf0;totalMemory[402] = 8'hf3;totalMemory[403] = 8'hec;totalMemory[404] = 8'he7;totalMemory[405] = 8'hbe;totalMemory[406] = 8'hb5;totalMemory[407] = 8'hb1;totalMemory[408] = 8'h6e;totalMemory[409] = 8'h65;totalMemory[410] = 8'h5d;totalMemory[411] = 8'h3d;totalMemory[412] = 8'h38;totalMemory[413] = 8'h2a;totalMemory[414] = 8'h39;totalMemory[415] = 8'h34;totalMemory[416] = 8'h16;totalMemory[417] = 8'h56;totalMemory[418] = 8'h4d;totalMemory[419] = 8'h17;totalMemory[420] = 8'h84;totalMemory[421] = 8'h73;totalMemory[422] = 8'h24;totalMemory[423] = 8'ha7;totalMemory[424] = 8'h8f;totalMemory[425] = 8'h25;totalMemory[426] = 8'hb8;totalMemory[427] = 8'h9b;totalMemory[428] = 8'h24;totalMemory[429] = 8'hb6;totalMemory[430] = 8'h9a;totalMemory[431] = 8'h22;totalMemory[432] = 8'ha6;totalMemory[433] = 8'h8c;totalMemory[434] = 8'h18;totalMemory[435] = 8'h95;totalMemory[436] = 8'h80;totalMemory[437] = 8'h11;totalMemory[438] = 8'h9a;totalMemory[439] = 8'h84;totalMemory[440] = 8'h10;totalMemory[441] = 8'hb1;totalMemory[442] = 8'h93;totalMemory[443] = 8'h14;totalMemory[444] = 8'hc1;totalMemory[445] = 8'h9d;totalMemory[446] = 8'h15;totalMemory[447] = 8'hc5;totalMemory[448] = 8'h9c;totalMemory[449] = 8'hf;totalMemory[450] = 8'hc6;totalMemory[451] = 8'h9a;totalMemory[452] = 8'h9;totalMemory[453] = 8'hce;totalMemory[454] = 8'ha0;totalMemory[455] = 8'hb;totalMemory[456] = 8'hdb;totalMemory[457] = 8'hab;totalMemory[458] = 8'h10;totalMemory[459] = 8'he5;totalMemory[460] = 8'hb4;totalMemory[461] = 8'he;totalMemory[462] = 8'he7;totalMemory[463] = 8'hb5;totalMemory[464] = 8'h6;totalMemory[465] = 8'he5;totalMemory[466] = 8'hb3;totalMemory[467] = 8'h1;totalMemory[468] = 8'he4;totalMemory[469] = 8'hb1;totalMemory[470] = 8'h0;totalMemory[471] = 8'he2;totalMemory[472] = 8'haf;totalMemory[473] = 8'h0;totalMemory[474] = 8'he0;totalMemory[475] = 8'haf;totalMemory[476] = 8'h0;totalMemory[477] = 8'hdd;totalMemory[478] = 8'hae;totalMemory[479] = 8'h0;totalMemory[480] = 8'hf3;totalMemory[481] = 8'hd1;totalMemory[482] = 8'hd4;totalMemory[483] = 8'hf6;totalMemory[484] = 8'hd2;totalMemory[485] = 8'hd3;totalMemory[486] = 8'hf8;totalMemory[487] = 8'hd5;totalMemory[488] = 8'hd5;totalMemory[489] = 8'hf9;totalMemory[490] = 8'hd8;totalMemory[491] = 8'hd7;totalMemory[492] = 8'hfc;totalMemory[493] = 8'hde;totalMemory[494] = 8'hdd;totalMemory[495] = 8'hfe;totalMemory[496] = 8'he9;totalMemory[497] = 8'he9;totalMemory[498] = 8'hff;totalMemory[499] = 8'hf1;totalMemory[500] = 8'hf1;totalMemory[501] = 8'hff;totalMemory[502] = 8'hef;totalMemory[503] = 8'hee;totalMemory[504] = 8'hff;totalMemory[505] = 8'hec;totalMemory[506] = 8'hea;totalMemory[507] = 8'hff;totalMemory[508] = 8'hee;totalMemory[509] = 8'hea;totalMemory[510] = 8'hff;totalMemory[511] = 8'hee;totalMemory[512] = 8'he9;totalMemory[513] = 8'hff;totalMemory[514] = 8'hf0;totalMemory[515] = 8'heb;totalMemory[516] = 8'hff;totalMemory[517] = 8'hf4;totalMemory[518] = 8'hf1;totalMemory[519] = 8'hef;totalMemory[520] = 8'he7;totalMemory[521] = 8'he4;totalMemory[522] = 8'hbc;totalMemory[523] = 8'hb2;totalMemory[524] = 8'hae;totalMemory[525] = 8'h72;totalMemory[526] = 8'h67;totalMemory[527] = 8'h62;totalMemory[528] = 8'h40;totalMemory[529] = 8'h38;totalMemory[530] = 8'h2d;totalMemory[531] = 8'h35;totalMemory[532] = 8'h31;totalMemory[533] = 8'h1b;totalMemory[534] = 8'h49;totalMemory[535] = 8'h42;totalMemory[536] = 8'h16;totalMemory[537] = 8'h79;totalMemory[538] = 8'h6a;totalMemory[539] = 8'h1f;totalMemory[540] = 8'ha6;totalMemory[541] = 8'h8f;totalMemory[542] = 8'h2a;totalMemory[543] = 8'hba;totalMemory[544] = 8'h9e;totalMemory[545] = 8'h27;totalMemory[546] = 8'hb9;totalMemory[547] = 8'h9d;totalMemory[548] = 8'h22;totalMemory[549] = 8'ha8;totalMemory[550] = 8'h91;totalMemory[551] = 8'h21;totalMemory[552] = 8'h95;totalMemory[553] = 8'h82;totalMemory[554] = 8'h16;totalMemory[555] = 8'h94;totalMemory[556] = 8'h82;totalMemory[557] = 8'h12;totalMemory[558] = 8'ha6;totalMemory[559] = 8'h8f;totalMemory[560] = 8'h19;totalMemory[561] = 8'hba;totalMemory[562] = 8'h9a;totalMemory[563] = 8'h1c;totalMemory[564] = 8'hc2;totalMemory[565] = 8'h9c;totalMemory[566] = 8'h17;totalMemory[567] = 8'hc5;totalMemory[568] = 8'h9b;totalMemory[569] = 8'h13;totalMemory[570] = 8'hcc;totalMemory[571] = 8'ha0;totalMemory[572] = 8'h12;totalMemory[573] = 8'hd6;totalMemory[574] = 8'ha7;totalMemory[575] = 8'h11;totalMemory[576] = 8'he1;totalMemory[577] = 8'hb1;totalMemory[578] = 8'hf;totalMemory[579] = 8'he8;totalMemory[580] = 8'hb7;totalMemory[581] = 8'ha;totalMemory[582] = 8'he7;totalMemory[583] = 8'hb4;totalMemory[584] = 8'h4;totalMemory[585] = 8'he4;totalMemory[586] = 8'hb0;totalMemory[587] = 8'h1;totalMemory[588] = 8'he1;totalMemory[589] = 8'hae;totalMemory[590] = 8'h0;totalMemory[591] = 8'hdf;totalMemory[592] = 8'had;totalMemory[593] = 8'h0;totalMemory[594] = 8'hdc;totalMemory[595] = 8'hac;totalMemory[596] = 8'h0;totalMemory[597] = 8'hd4;totalMemory[598] = 8'ha9;totalMemory[599] = 8'h1;totalMemory[600] = 8'hff;totalMemory[601] = 8'he6;totalMemory[602] = 8'he8;totalMemory[603] = 8'hff;totalMemory[604] = 8'he1;totalMemory[605] = 8'he1;totalMemory[606] = 8'hff;totalMemory[607] = 8'he6;totalMemory[608] = 8'he5;totalMemory[609] = 8'hff;totalMemory[610] = 8'hec;totalMemory[611] = 8'hea;totalMemory[612] = 8'hff;totalMemory[613] = 8'hee;totalMemory[614] = 8'hec;totalMemory[615] = 8'hff;totalMemory[616] = 8'hf3;totalMemory[617] = 8'hf1;totalMemory[618] = 8'hff;totalMemory[619] = 8'hf5;totalMemory[620] = 8'hf3;totalMemory[621] = 8'hff;totalMemory[622] = 8'hf0;totalMemory[623] = 8'hed;totalMemory[624] = 8'hff;totalMemory[625] = 8'hee;totalMemory[626] = 8'heb;totalMemory[627] = 8'hff;totalMemory[628] = 8'hf2;totalMemory[629] = 8'hee;totalMemory[630] = 8'hff;totalMemory[631] = 8'hf6;totalMemory[632] = 8'hf3;totalMemory[633] = 8'hff;totalMemory[634] = 8'hf7;totalMemory[635] = 8'hf4;totalMemory[636] = 8'heb;totalMemory[637] = 8'he0;totalMemory[638] = 8'hdd;totalMemory[639] = 8'hb0;totalMemory[640] = 8'ha3;totalMemory[641] = 8'h9f;totalMemory[642] = 8'h69;totalMemory[643] = 8'h5d;totalMemory[644] = 8'h58;totalMemory[645] = 8'h3d;totalMemory[646] = 8'h34;totalMemory[647] = 8'h2c;totalMemory[648] = 8'h33;totalMemory[649] = 8'h2d;totalMemory[650] = 8'h1b;totalMemory[651] = 8'h3f;totalMemory[652] = 8'h39;totalMemory[653] = 8'h17;totalMemory[654] = 8'h68;totalMemory[655] = 8'h5c;totalMemory[656] = 8'h21;totalMemory[657] = 8'ha1;totalMemory[658] = 8'h8b;totalMemory[659] = 8'h30;totalMemory[660] = 8'hc1;totalMemory[661] = 8'ha4;totalMemory[662] = 8'h34;totalMemory[663] = 8'hbe;totalMemory[664] = 8'h9f;totalMemory[665] = 8'h28;totalMemory[666] = 8'ha9;totalMemory[667] = 8'h8f;totalMemory[668] = 8'h1b;totalMemory[669] = 8'h93;totalMemory[670] = 8'h80;totalMemory[671] = 8'h17;totalMemory[672] = 8'h8d;totalMemory[673] = 8'h7d;totalMemory[674] = 8'h16;totalMemory[675] = 8'h9b;totalMemory[676] = 8'h89;totalMemory[677] = 8'h1b;totalMemory[678] = 8'hb1;totalMemory[679] = 8'h98;totalMemory[680] = 8'h22;totalMemory[681] = 8'hbd;totalMemory[682] = 8'h9c;totalMemory[683] = 8'h1f;totalMemory[684] = 8'hc3;totalMemory[685] = 8'h9a;totalMemory[686] = 8'h19;totalMemory[687] = 8'hcc;totalMemory[688] = 8'ha1;totalMemory[689] = 8'h1a;totalMemory[690] = 8'hd7;totalMemory[691] = 8'haa;totalMemory[692] = 8'h1c;totalMemory[693] = 8'hdb;totalMemory[694] = 8'hac;totalMemory[695] = 8'h15;totalMemory[696] = 8'hde;totalMemory[697] = 8'had;totalMemory[698] = 8'hc;totalMemory[699] = 8'hdf;totalMemory[700] = 8'hae;totalMemory[701] = 8'h5;totalMemory[702] = 8'hdd;totalMemory[703] = 8'hab;totalMemory[704] = 8'h1;totalMemory[705] = 8'hde;totalMemory[706] = 8'hab;totalMemory[707] = 8'h0;totalMemory[708] = 8'hde;totalMemory[709] = 8'hac;totalMemory[710] = 8'h0;totalMemory[711] = 8'hdc;totalMemory[712] = 8'hab;totalMemory[713] = 8'h0;totalMemory[714] = 8'hd4;totalMemory[715] = 8'ha8;totalMemory[716] = 8'h1;totalMemory[717] = 8'hc7;totalMemory[718] = 8'ha1;totalMemory[719] = 8'h3;totalMemory[720] = 8'hfe;totalMemory[721] = 8'he7;totalMemory[722] = 8'he8;totalMemory[723] = 8'hff;totalMemory[724] = 8'he2;totalMemory[725] = 8'he3;totalMemory[726] = 8'hff;totalMemory[727] = 8'he9;totalMemory[728] = 8'hea;totalMemory[729] = 8'hff;totalMemory[730] = 8'hec;totalMemory[731] = 8'hec;totalMemory[732] = 8'hff;totalMemory[733] = 8'hf1;totalMemory[734] = 8'hef;totalMemory[735] = 8'hff;totalMemory[736] = 8'hf5;totalMemory[737] = 8'hf3;totalMemory[738] = 8'hff;totalMemory[739] = 8'hf1;totalMemory[740] = 8'hee;totalMemory[741] = 8'hff;totalMemory[742] = 8'heb;totalMemory[743] = 8'he8;totalMemory[744] = 8'hff;totalMemory[745] = 8'hec;totalMemory[746] = 8'he8;totalMemory[747] = 8'hff;totalMemory[748] = 8'hf2;totalMemory[749] = 8'hee;totalMemory[750] = 8'hf9;totalMemory[751] = 8'hef;totalMemory[752] = 8'hed;totalMemory[753] = 8'hdc;totalMemory[754] = 8'hd2;totalMemory[755] = 8'hcf;totalMemory[756] = 8'ha0;totalMemory[757] = 8'h95;totalMemory[758] = 8'h90;totalMemory[759] = 8'h5c;totalMemory[760] = 8'h52;totalMemory[761] = 8'h4b;totalMemory[762] = 8'h39;totalMemory[763] = 8'h32;totalMemory[764] = 8'h28;totalMemory[765] = 8'h33;totalMemory[766] = 8'h2e;totalMemory[767] = 8'h20;totalMemory[768] = 8'h3b;totalMemory[769] = 8'h35;totalMemory[770] = 8'h1a;totalMemory[771] = 8'h5c;totalMemory[772] = 8'h51;totalMemory[773] = 8'h1f;totalMemory[774] = 8'h96;totalMemory[775] = 8'h83;totalMemory[776] = 8'h37;totalMemory[777] = 8'hc3;totalMemory[778] = 8'ha5;totalMemory[779] = 8'h3f;totalMemory[780] = 8'hc6;totalMemory[781] = 8'ha5;totalMemory[782] = 8'h36;totalMemory[783] = 8'hae;totalMemory[784] = 8'h90;totalMemory[785] = 8'h28;totalMemory[786] = 8'h92;totalMemory[787] = 8'h7a;totalMemory[788] = 8'h18;totalMemory[789] = 8'h88;totalMemory[790] = 8'h77;totalMemory[791] = 8'h17;totalMemory[792] = 8'h94;totalMemory[793] = 8'h83;totalMemory[794] = 8'h1e;totalMemory[795] = 8'ha7;totalMemory[796] = 8'h91;totalMemory[797] = 8'h22;totalMemory[798] = 8'hb4;totalMemory[799] = 8'h97;totalMemory[800] = 8'h21;totalMemory[801] = 8'hbb;totalMemory[802] = 8'h99;totalMemory[803] = 8'h1e;totalMemory[804] = 8'hc6;totalMemory[805] = 8'h9e;totalMemory[806] = 8'h1e;totalMemory[807] = 8'hd4;totalMemory[808] = 8'ha8;totalMemory[809] = 8'h1e;totalMemory[810] = 8'hdd;totalMemory[811] = 8'haf;totalMemory[812] = 8'h1d;totalMemory[813] = 8'hdc;totalMemory[814] = 8'hac;totalMemory[815] = 8'h14;totalMemory[816] = 8'hd7;totalMemory[817] = 8'ha7;totalMemory[818] = 8'ha;totalMemory[819] = 8'hd3;totalMemory[820] = 8'ha3;totalMemory[821] = 8'h4;totalMemory[822] = 8'hd0;totalMemory[823] = 8'ha3;totalMemory[824] = 8'h1;totalMemory[825] = 8'hd5;totalMemory[826] = 8'ha6;totalMemory[827] = 8'h2;totalMemory[828] = 8'hd4;totalMemory[829] = 8'ha6;totalMemory[830] = 8'h2;totalMemory[831] = 8'hce;totalMemory[832] = 8'ha1;totalMemory[833] = 8'h0;totalMemory[834] = 8'hc4;totalMemory[835] = 8'h9e;totalMemory[836] = 8'h3;totalMemory[837] = 8'hb7;totalMemory[838] = 8'h9a;totalMemory[839] = 8'h8;totalMemory[840] = 8'hf8;totalMemory[841] = 8'hda;totalMemory[842] = 8'hdc;totalMemory[843] = 8'hfb;totalMemory[844] = 8'hdd;totalMemory[845] = 8'hdf;totalMemory[846] = 8'hfe;totalMemory[847] = 8'he5;totalMemory[848] = 8'he8;totalMemory[849] = 8'hff;totalMemory[850] = 8'he7;totalMemory[851] = 8'he8;totalMemory[852] = 8'hff;totalMemory[853] = 8'hea;totalMemory[854] = 8'hea;totalMemory[855] = 8'hff;totalMemory[856] = 8'hee;totalMemory[857] = 8'hec;totalMemory[858] = 8'hff;totalMemory[859] = 8'hec;totalMemory[860] = 8'hea;totalMemory[861] = 8'hff;totalMemory[862] = 8'heb;totalMemory[863] = 8'he9;totalMemory[864] = 8'hfe;totalMemory[865] = 8'hec;totalMemory[866] = 8'hea;totalMemory[867] = 8'hed;totalMemory[868] = 8'hde;totalMemory[869] = 8'hdb;totalMemory[870] = 8'hc3;totalMemory[871] = 8'hb5;totalMemory[872] = 8'hb1;totalMemory[873] = 8'h85;totalMemory[874] = 8'h79;totalMemory[875] = 8'h72;totalMemory[876] = 8'h4e;totalMemory[877] = 8'h45;totalMemory[878] = 8'h3c;totalMemory[879] = 8'h36;totalMemory[880] = 8'h31;totalMemory[881] = 8'h25;totalMemory[882] = 8'h33;totalMemory[883] = 8'h30;totalMemory[884] = 8'h20;totalMemory[885] = 8'h37;totalMemory[886] = 8'h32;totalMemory[887] = 8'h1f;totalMemory[888] = 8'h54;totalMemory[889] = 8'h4b;totalMemory[890] = 8'h2b;totalMemory[891] = 8'h94;totalMemory[892] = 8'h85;totalMemory[893] = 8'h4e;totalMemory[894] = 8'hc8;totalMemory[895] = 8'hb1;totalMemory[896] = 8'h62;totalMemory[897] = 8'hd0;totalMemory[898] = 8'haf;totalMemory[899] = 8'h4d;totalMemory[900] = 8'hbb;totalMemory[901] = 8'h98;totalMemory[902] = 8'h33;totalMemory[903] = 8'h99;totalMemory[904] = 8'h7d;totalMemory[905] = 8'h22;totalMemory[906] = 8'h87;totalMemory[907] = 8'h72;totalMemory[908] = 8'h1b;totalMemory[909] = 8'h92;totalMemory[910] = 8'h7f;totalMemory[911] = 8'h22;totalMemory[912] = 8'ha3;totalMemory[913] = 8'h8f;totalMemory[914] = 8'h2a;totalMemory[915] = 8'hb0;totalMemory[916] = 8'h96;totalMemory[917] = 8'h28;totalMemory[918] = 8'hb9;totalMemory[919] = 8'h98;totalMemory[920] = 8'h23;totalMemory[921] = 8'hc2;totalMemory[922] = 8'h9e;totalMemory[923] = 8'h24;totalMemory[924] = 8'hcc;totalMemory[925] = 8'ha5;totalMemory[926] = 8'h25;totalMemory[927] = 8'hd4;totalMemory[928] = 8'hab;totalMemory[929] = 8'h21;totalMemory[930] = 8'hd7;totalMemory[931] = 8'had;totalMemory[932] = 8'h1d;totalMemory[933] = 8'hd2;totalMemory[934] = 8'ha7;totalMemory[935] = 8'h17;totalMemory[936] = 8'hc9;totalMemory[937] = 8'h9f;totalMemory[938] = 8'hd;totalMemory[939] = 8'hc4;totalMemory[940] = 8'h9a;totalMemory[941] = 8'h6;totalMemory[942] = 8'hc4;totalMemory[943] = 8'h9a;totalMemory[944] = 8'h3;totalMemory[945] = 8'hc8;totalMemory[946] = 8'h9e;totalMemory[947] = 8'h3;totalMemory[948] = 8'hc6;totalMemory[949] = 8'h9e;totalMemory[950] = 8'h2;totalMemory[951] = 8'hc1;totalMemory[952] = 8'h9b;totalMemory[953] = 8'h2;totalMemory[954] = 8'hb9;totalMemory[955] = 8'h9a;totalMemory[956] = 8'h7;totalMemory[957] = 8'hac;totalMemory[958] = 8'h98;totalMemory[959] = 8'h10;totalMemory[960] = 8'hf6;totalMemory[961] = 8'hd8;totalMemory[962] = 8'hda;totalMemory[963] = 8'hfa;totalMemory[964] = 8'hdb;totalMemory[965] = 8'hdd;totalMemory[966] = 8'hfe;totalMemory[967] = 8'he1;totalMemory[968] = 8'he2;totalMemory[969] = 8'hfe;totalMemory[970] = 8'he3;totalMemory[971] = 8'he2;totalMemory[972] = 8'hfc;totalMemory[973] = 8'he2;totalMemory[974] = 8'he0;totalMemory[975] = 8'hfd;totalMemory[976] = 8'he5;totalMemory[977] = 8'he3;totalMemory[978] = 8'hff;totalMemory[979] = 8'hea;totalMemory[980] = 8'he9;totalMemory[981] = 8'hfb;totalMemory[982] = 8'heb;totalMemory[983] = 8'hea;totalMemory[984] = 8'hde;totalMemory[985] = 8'hcd;totalMemory[986] = 8'hcd;totalMemory[987] = 8'ha3;totalMemory[988] = 8'h93;totalMemory[989] = 8'h8f;totalMemory[990] = 8'h67;totalMemory[991] = 8'h5b;totalMemory[992] = 8'h54;totalMemory[993] = 8'h42;totalMemory[994] = 8'h3c;totalMemory[995] = 8'h31;totalMemory[996] = 8'h36;totalMemory[997] = 8'h32;totalMemory[998] = 8'h25;totalMemory[999] = 8'h37;totalMemory[1000] = 8'h35;totalMemory[1001] = 8'h24;totalMemory[1002] = 8'h3a;totalMemory[1003] = 8'h36;totalMemory[1004] = 8'h21;totalMemory[1005] = 8'h4a;totalMemory[1006] = 8'h43;totalMemory[1007] = 8'h2b;totalMemory[1008] = 8'h89;totalMemory[1009] = 8'h7b;totalMemory[1010] = 8'h5b;totalMemory[1011] = 8'hd2;totalMemory[1012] = 8'hbd;totalMemory[1013] = 8'h8e;totalMemory[1014] = 8'he2;totalMemory[1015] = 8'hc8;totalMemory[1016] = 8'h89;totalMemory[1017] = 8'hc7;totalMemory[1018] = 8'ha7;totalMemory[1019] = 8'h59;totalMemory[1020] = 8'ha4;totalMemory[1021] = 8'h85;totalMemory[1022] = 8'h32;totalMemory[1023] = 8'h8b;totalMemory[1024] = 8'h72;totalMemory[1025] = 8'h23;totalMemory[1026] = 8'h90;totalMemory[1027] = 8'h7a;totalMemory[1028] = 8'h28;totalMemory[1029] = 8'ha5;totalMemory[1030] = 8'h8e;totalMemory[1031] = 8'h2e;totalMemory[1032] = 8'hb3;totalMemory[1033] = 8'h99;totalMemory[1034] = 8'h2e;totalMemory[1035] = 8'hbc;totalMemory[1036] = 8'h9e;totalMemory[1037] = 8'h2e;totalMemory[1038] = 8'hc3;totalMemory[1039] = 8'ha1;totalMemory[1040] = 8'h2d;totalMemory[1041] = 8'hcb;totalMemory[1042] = 8'ha6;totalMemory[1043] = 8'h2b;totalMemory[1044] = 8'hcf;totalMemory[1045] = 8'ha9;totalMemory[1046] = 8'h29;totalMemory[1047] = 8'hcc;totalMemory[1048] = 8'ha8;totalMemory[1049] = 8'h23;totalMemory[1050] = 8'hc3;totalMemory[1051] = 8'ha1;totalMemory[1052] = 8'h1b;totalMemory[1053] = 8'hb4;totalMemory[1054] = 8'h95;totalMemory[1055] = 8'h14;totalMemory[1056] = 8'hac;totalMemory[1057] = 8'h8e;totalMemory[1058] = 8'he;totalMemory[1059] = 8'hb0;totalMemory[1060] = 8'h8f;totalMemory[1061] = 8'hb;totalMemory[1062] = 8'hb7;totalMemory[1063] = 8'h93;totalMemory[1064] = 8'h8;totalMemory[1065] = 8'hbe;totalMemory[1066] = 8'h97;totalMemory[1067] = 8'h5;totalMemory[1068] = 8'hc2;totalMemory[1069] = 8'h9c;totalMemory[1070] = 8'h6;totalMemory[1071] = 8'hc0;totalMemory[1072] = 8'h9f;totalMemory[1073] = 8'h8;totalMemory[1074] = 8'hb4;totalMemory[1075] = 8'h9c;totalMemory[1076] = 8'hc;totalMemory[1077] = 8'ha1;totalMemory[1078] = 8'h98;totalMemory[1079] = 8'h15;totalMemory[1080] = 8'hf5;totalMemory[1081] = 8'hda;totalMemory[1082] = 8'hda;totalMemory[1083] = 8'hfa;totalMemory[1084] = 8'hde;totalMemory[1085] = 8'hde;totalMemory[1086] = 8'hf6;totalMemory[1087] = 8'hdb;totalMemory[1088] = 8'hd9;totalMemory[1089] = 8'hed;totalMemory[1090] = 8'hd3;totalMemory[1091] = 8'hd0;totalMemory[1092] = 8'hee;totalMemory[1093] = 8'hd7;totalMemory[1094] = 8'hd3;totalMemory[1095] = 8'hf7;totalMemory[1096] = 8'he2;totalMemory[1097] = 8'hde;totalMemory[1098] = 8'hf0;totalMemory[1099] = 8'he1;totalMemory[1100] = 8'hde;totalMemory[1101] = 8'hcc;totalMemory[1102] = 8'hbf;totalMemory[1103] = 8'hbd;totalMemory[1104] = 8'h8a;totalMemory[1105] = 8'h7d;totalMemory[1106] = 8'h7a;totalMemory[1107] = 8'h4f;totalMemory[1108] = 8'h45;totalMemory[1109] = 8'h3e;totalMemory[1110] = 8'h3a;totalMemory[1111] = 8'h33;totalMemory[1112] = 8'h29;totalMemory[1113] = 8'h38;totalMemory[1114] = 8'h35;totalMemory[1115] = 8'h28;totalMemory[1116] = 8'h3a;totalMemory[1117] = 8'h37;totalMemory[1118] = 8'h27;totalMemory[1119] = 8'h40;totalMemory[1120] = 8'h3b;totalMemory[1121] = 8'h28;totalMemory[1122] = 8'h56;totalMemory[1123] = 8'h4d;totalMemory[1124] = 8'h38;totalMemory[1125] = 8'h85;totalMemory[1126] = 8'h78;totalMemory[1127] = 8'h61;totalMemory[1128] = 8'hc4;totalMemory[1129] = 8'hb1;totalMemory[1130] = 8'h94;totalMemory[1131] = 8'he7;totalMemory[1132] = 8'hcf;totalMemory[1133] = 8'ha7;totalMemory[1134] = 8'hd7;totalMemory[1135] = 8'hba;totalMemory[1136] = 8'h87;totalMemory[1137] = 8'hb0;totalMemory[1138] = 8'h91;totalMemory[1139] = 8'h52;totalMemory[1140] = 8'h93;totalMemory[1141] = 8'h75;totalMemory[1142] = 8'h2e;totalMemory[1143] = 8'h8f;totalMemory[1144] = 8'h75;totalMemory[1145] = 8'h2d;totalMemory[1146] = 8'ha0;totalMemory[1147] = 8'h88;totalMemory[1148] = 8'h38;totalMemory[1149] = 8'hb1;totalMemory[1150] = 8'h96;totalMemory[1151] = 8'h39;totalMemory[1152] = 8'hbc;totalMemory[1153] = 8'h9f;totalMemory[1154] = 8'h37;totalMemory[1155] = 8'hc4;totalMemory[1156] = 8'ha5;totalMemory[1157] = 8'h3a;totalMemory[1158] = 8'hc6;totalMemory[1159] = 8'ha5;totalMemory[1160] = 8'h37;totalMemory[1161] = 8'hc3;totalMemory[1162] = 8'ha2;totalMemory[1163] = 8'h2e;totalMemory[1164] = 8'hbd;totalMemory[1165] = 8'h9e;totalMemory[1166] = 8'h26;totalMemory[1167] = 8'hae;totalMemory[1168] = 8'h94;totalMemory[1169] = 8'h1b;totalMemory[1170] = 8'h9c;totalMemory[1171] = 8'h85;totalMemory[1172] = 8'he;totalMemory[1173] = 8'h90;totalMemory[1174] = 8'h7b;totalMemory[1175] = 8'h8;totalMemory[1176] = 8'h95;totalMemory[1177] = 8'h7f;totalMemory[1178] = 8'ha;totalMemory[1179] = 8'ha6;totalMemory[1180] = 8'h8b;totalMemory[1181] = 8'he;totalMemory[1182] = 8'hb5;totalMemory[1183] = 8'h95;totalMemory[1184] = 8'he;totalMemory[1185] = 8'hbf;totalMemory[1186] = 8'h9c;totalMemory[1187] = 8'hc;totalMemory[1188] = 8'hc1;totalMemory[1189] = 8'ha0;totalMemory[1190] = 8'hc;totalMemory[1191] = 8'hbb;totalMemory[1192] = 8'ha0;totalMemory[1193] = 8'he;totalMemory[1194] = 8'ha9;totalMemory[1195] = 8'h9b;totalMemory[1196] = 8'h12;totalMemory[1197] = 8'h90;totalMemory[1198] = 8'h91;totalMemory[1199] = 8'h19;totalMemory[1200] = 8'hcc;totalMemory[1201] = 8'hb9;totalMemory[1202] = 8'hb4;totalMemory[1203] = 8'hc5;totalMemory[1204] = 8'hb2;totalMemory[1205] = 8'had;totalMemory[1206] = 8'hb7;totalMemory[1207] = 8'ha4;totalMemory[1208] = 8'h9e;totalMemory[1209] = 8'hb9;totalMemory[1210] = 8'ha8;totalMemory[1211] = 8'ha0;totalMemory[1212] = 8'hc5;totalMemory[1213] = 8'hb6;totalMemory[1214] = 8'hae;totalMemory[1215] = 8'hc3;totalMemory[1216] = 8'hb6;totalMemory[1217] = 8'had;totalMemory[1218] = 8'ha5;totalMemory[1219] = 8'h98;totalMemory[1220] = 8'h91;totalMemory[1221] = 8'h6f;totalMemory[1222] = 8'h65;totalMemory[1223] = 8'h5e;totalMemory[1224] = 8'h43;totalMemory[1225] = 8'h3b;totalMemory[1226] = 8'h34;totalMemory[1227] = 8'h37;totalMemory[1228] = 8'h31;totalMemory[1229] = 8'h27;totalMemory[1230] = 8'h3b;totalMemory[1231] = 8'h36;totalMemory[1232] = 8'h29;totalMemory[1233] = 8'h3b;totalMemory[1234] = 8'h37;totalMemory[1235] = 8'h28;totalMemory[1236] = 8'h41;totalMemory[1237] = 8'h3c;totalMemory[1238] = 8'h2a;totalMemory[1239] = 8'h60;totalMemory[1240] = 8'h56;totalMemory[1241] = 8'h43;totalMemory[1242] = 8'h9b;totalMemory[1243] = 8'h8b;totalMemory[1244] = 8'h79;totalMemory[1245] = 8'hd0;totalMemory[1246] = 8'hbc;totalMemory[1247] = 8'had;totalMemory[1248] = 8'he8;totalMemory[1249] = 8'hce;totalMemory[1250] = 8'hba;totalMemory[1251] = 8'hde;totalMemory[1252] = 8'hc1;totalMemory[1253] = 8'ha0;totalMemory[1254] = 8'hbc;totalMemory[1255] = 8'h9e;totalMemory[1256] = 8'h71;totalMemory[1257] = 8'h9b;totalMemory[1258] = 8'h7e;totalMemory[1259] = 8'h45;totalMemory[1260] = 8'h91;totalMemory[1261] = 8'h76;totalMemory[1262] = 8'h34;totalMemory[1263] = 8'h9f;totalMemory[1264] = 8'h83;totalMemory[1265] = 8'h3b;totalMemory[1266] = 8'haf;totalMemory[1267] = 8'h93;totalMemory[1268] = 8'h44;totalMemory[1269] = 8'hb9;totalMemory[1270] = 8'h9d;totalMemory[1271] = 8'h45;totalMemory[1272] = 8'hbf;totalMemory[1273] = 8'ha2;totalMemory[1274] = 8'h45;totalMemory[1275] = 8'hbd;totalMemory[1276] = 8'ha0;totalMemory[1277] = 8'h42;totalMemory[1278] = 8'hb1;totalMemory[1279] = 8'h96;totalMemory[1280] = 8'h36;totalMemory[1281] = 8'ha0;totalMemory[1282] = 8'h89;totalMemory[1283] = 8'h27;totalMemory[1284] = 8'h90;totalMemory[1285] = 8'h7e;totalMemory[1286] = 8'h1c;totalMemory[1287] = 8'h82;totalMemory[1288] = 8'h76;totalMemory[1289] = 8'h14;totalMemory[1290] = 8'h7b;totalMemory[1291] = 8'h72;totalMemory[1292] = 8'he;totalMemory[1293] = 8'h81;totalMemory[1294] = 8'h76;totalMemory[1295] = 8'he;totalMemory[1296] = 8'h95;totalMemory[1297] = 8'h83;totalMemory[1298] = 8'h11;totalMemory[1299] = 8'had;totalMemory[1300] = 8'h94;totalMemory[1301] = 8'h12;totalMemory[1302] = 8'hbd;totalMemory[1303] = 8'h9e;totalMemory[1304] = 8'h11;totalMemory[1305] = 8'hc4;totalMemory[1306] = 8'ha1;totalMemory[1307] = 8'hd;totalMemory[1308] = 8'hbe;totalMemory[1309] = 8'ha0;totalMemory[1310] = 8'he;totalMemory[1311] = 8'hac;totalMemory[1312] = 8'h9b;totalMemory[1313] = 8'h12;totalMemory[1314] = 8'h95;totalMemory[1315] = 8'h92;totalMemory[1316] = 8'h17;totalMemory[1317] = 8'h7b;totalMemory[1318] = 8'h87;totalMemory[1319] = 8'h1c;totalMemory[1320] = 8'h7c;totalMemory[1321] = 8'h71;totalMemory[1322] = 8'h68;totalMemory[1323] = 8'h69;totalMemory[1324] = 8'h5e;totalMemory[1325] = 8'h53;totalMemory[1326] = 8'h61;totalMemory[1327] = 8'h56;totalMemory[1328] = 8'h4a;totalMemory[1329] = 8'h6f;totalMemory[1330] = 8'h64;totalMemory[1331] = 8'h59;totalMemory[1332] = 8'h74;totalMemory[1333] = 8'h6a;totalMemory[1334] = 8'h5f;totalMemory[1335] = 8'h63;totalMemory[1336] = 8'h5b;totalMemory[1337] = 8'h4f;totalMemory[1338] = 8'h4c;totalMemory[1339] = 8'h44;totalMemory[1340] = 8'h38;totalMemory[1341] = 8'h38;totalMemory[1342] = 8'h30;totalMemory[1343] = 8'h26;totalMemory[1344] = 8'h35;totalMemory[1345] = 8'h2e;totalMemory[1346] = 8'h22;totalMemory[1347] = 8'h3b;totalMemory[1348] = 8'h34;totalMemory[1349] = 8'h27;totalMemory[1350] = 8'h3f;totalMemory[1351] = 8'h38;totalMemory[1352] = 8'h2a;totalMemory[1353] = 8'h49;totalMemory[1354] = 8'h41;totalMemory[1355] = 8'h32;totalMemory[1356] = 8'h69;totalMemory[1357] = 8'h5e;totalMemory[1358] = 8'h4d;totalMemory[1359] = 8'ha0;totalMemory[1360] = 8'h8f;totalMemory[1361] = 8'h7f;totalMemory[1362] = 8'hda;totalMemory[1363] = 8'hc5;totalMemory[1364] = 8'hb7;totalMemory[1365] = 8'hf7;totalMemory[1366] = 8'hdf;totalMemory[1367] = 8'hd5;totalMemory[1368] = 8'hf5;totalMemory[1369] = 8'hda;totalMemory[1370] = 8'hcb;totalMemory[1371] = 8'hd4;totalMemory[1372] = 8'hb6;totalMemory[1373] = 8'h9b;totalMemory[1374] = 8'ha5;totalMemory[1375] = 8'h88;totalMemory[1376] = 8'h60;totalMemory[1377] = 8'h92;totalMemory[1378] = 8'h77;totalMemory[1379] = 8'h43;totalMemory[1380] = 8'ha0;totalMemory[1381] = 8'h86;totalMemory[1382] = 8'h4a;totalMemory[1383] = 8'hb6;totalMemory[1384] = 8'h9d;totalMemory[1385] = 8'h5a;totalMemory[1386] = 8'hc1;totalMemory[1387] = 8'ha8;totalMemory[1388] = 8'h60;totalMemory[1389] = 8'hbb;totalMemory[1390] = 8'ha1;totalMemory[1391] = 8'h57;totalMemory[1392] = 8'ha8;totalMemory[1393] = 8'h8f;totalMemory[1394] = 8'h43;totalMemory[1395] = 8'h96;totalMemory[1396] = 8'h7f;totalMemory[1397] = 8'h31;totalMemory[1398] = 8'h88;totalMemory[1399] = 8'h74;totalMemory[1400] = 8'h25;totalMemory[1401] = 8'h79;totalMemory[1402] = 8'h6b;totalMemory[1403] = 8'h1a;totalMemory[1404] = 8'h6e;totalMemory[1405] = 8'h65;totalMemory[1406] = 8'h12;totalMemory[1407] = 8'h6e;totalMemory[1408] = 8'h6a;totalMemory[1409] = 8'h13;totalMemory[1410] = 8'h79;totalMemory[1411] = 8'h75;totalMemory[1412] = 8'h17;totalMemory[1413] = 8'h8c;totalMemory[1414] = 8'h83;totalMemory[1415] = 8'h1b;totalMemory[1416] = 8'ha3;totalMemory[1417] = 8'h92;totalMemory[1418] = 8'h1b;totalMemory[1419] = 8'hb6;totalMemory[1420] = 8'h9d;totalMemory[1421] = 8'h16;totalMemory[1422] = 8'hbe;totalMemory[1423] = 8'ha1;totalMemory[1424] = 8'h11;totalMemory[1425] = 8'hbd;totalMemory[1426] = 8'h9f;totalMemory[1427] = 8'he;totalMemory[1428] = 8'haf;totalMemory[1429] = 8'h99;totalMemory[1430] = 8'he;totalMemory[1431] = 8'h98;totalMemory[1432] = 8'h91;totalMemory[1433] = 8'h14;totalMemory[1434] = 8'h82;totalMemory[1435] = 8'h8a;totalMemory[1436] = 8'h1c;totalMemory[1437] = 8'h6d;totalMemory[1438] = 8'h82;totalMemory[1439] = 8'h23;totalMemory[1440] = 8'h40;totalMemory[1441] = 8'h3a;totalMemory[1442] = 8'h2e;totalMemory[1443] = 8'h3b;totalMemory[1444] = 8'h36;totalMemory[1445] = 8'h29;totalMemory[1446] = 8'h39;totalMemory[1447] = 8'h34;totalMemory[1448] = 8'h26;totalMemory[1449] = 8'h38;totalMemory[1450] = 8'h33;totalMemory[1451] = 8'h26;totalMemory[1452] = 8'h35;totalMemory[1453] = 8'h30;totalMemory[1454] = 8'h22;totalMemory[1455] = 8'h34;totalMemory[1456] = 8'h2d;totalMemory[1457] = 8'h1f;totalMemory[1458] = 8'h34;totalMemory[1459] = 8'h2d;totalMemory[1460] = 8'h1d;totalMemory[1461] = 8'h37;totalMemory[1462] = 8'h30;totalMemory[1463] = 8'h21;totalMemory[1464] = 8'h44;totalMemory[1465] = 8'h3a;totalMemory[1466] = 8'h2c;totalMemory[1467] = 8'h52;totalMemory[1468] = 8'h46;totalMemory[1469] = 8'h37;totalMemory[1470] = 8'h69;totalMemory[1471] = 8'h5b;totalMemory[1472] = 8'h4c;totalMemory[1473] = 8'h8c;totalMemory[1474] = 8'h7c;totalMemory[1475] = 8'h6f;totalMemory[1476] = 8'hb0;totalMemory[1477] = 8'h9e;totalMemory[1478] = 8'h92;totalMemory[1479] = 8'hd6;totalMemory[1480] = 8'hc0;totalMemory[1481] = 8'hb6;totalMemory[1482] = 8'hf3;totalMemory[1483] = 8'hdd;totalMemory[1484] = 8'hd4;totalMemory[1485] = 8'hfe;totalMemory[1486] = 8'he9;totalMemory[1487] = 8'he0;totalMemory[1488] = 8'hf1;totalMemory[1489] = 8'hd8;totalMemory[1490] = 8'hca;totalMemory[1491] = 8'hc2;totalMemory[1492] = 8'ha6;totalMemory[1493] = 8'h8d;totalMemory[1494] = 8'h9e;totalMemory[1495] = 8'h81;totalMemory[1496] = 8'h5d;totalMemory[1497] = 8'ha5;totalMemory[1498] = 8'h89;totalMemory[1499] = 8'h59;totalMemory[1500] = 8'hbb;totalMemory[1501] = 8'ha2;totalMemory[1502] = 8'h6d;totalMemory[1503] = 8'hc8;totalMemory[1504] = 8'hb4;totalMemory[1505] = 8'h7e;totalMemory[1506] = 8'hbf;totalMemory[1507] = 8'had;totalMemory[1508] = 8'h79;totalMemory[1509] = 8'h9a;totalMemory[1510] = 8'h8a;totalMemory[1511] = 8'h55;totalMemory[1512] = 8'h74;totalMemory[1513] = 8'h66;totalMemory[1514] = 8'h30;totalMemory[1515] = 8'h66;totalMemory[1516] = 8'h58;totalMemory[1517] = 8'h22;totalMemory[1518] = 8'h63;totalMemory[1519] = 8'h59;totalMemory[1520] = 8'h1e;totalMemory[1521] = 8'h61;totalMemory[1522] = 8'h5d;totalMemory[1523] = 8'h1b;totalMemory[1524] = 8'h66;totalMemory[1525] = 8'h64;totalMemory[1526] = 8'h19;totalMemory[1527] = 8'h76;totalMemory[1528] = 8'h73;totalMemory[1529] = 8'h19;totalMemory[1530] = 8'h8c;totalMemory[1531] = 8'h84;totalMemory[1532] = 8'h1d;totalMemory[1533] = 8'h9f;totalMemory[1534] = 8'h91;totalMemory[1535] = 8'h1e;totalMemory[1536] = 8'haa;totalMemory[1537] = 8'h97;totalMemory[1538] = 8'h16;totalMemory[1539] = 8'hb0;totalMemory[1540] = 8'h98;totalMemory[1541] = 8'hc;totalMemory[1542] = 8'hb3;totalMemory[1543] = 8'h9a;totalMemory[1544] = 8'hc;totalMemory[1545] = 8'had;totalMemory[1546] = 8'h97;totalMemory[1547] = 8'hf;totalMemory[1548] = 8'h9a;totalMemory[1549] = 8'h8f;totalMemory[1550] = 8'h12;totalMemory[1551] = 8'h83;totalMemory[1552] = 8'h89;totalMemory[1553] = 8'h1b;totalMemory[1554] = 8'h73;totalMemory[1555] = 8'h87;totalMemory[1556] = 8'h26;totalMemory[1557] = 8'h65;totalMemory[1558] = 8'h82;totalMemory[1559] = 8'h2c;totalMemory[1560] = 8'h36;totalMemory[1561] = 8'h34;totalMemory[1562] = 8'h26;totalMemory[1563] = 8'h36;totalMemory[1564] = 8'h35;totalMemory[1565] = 8'h26;totalMemory[1566] = 8'h2e;totalMemory[1567] = 8'h2c;totalMemory[1568] = 8'h1e;totalMemory[1569] = 8'h2b;totalMemory[1570] = 8'h27;totalMemory[1571] = 8'h18;totalMemory[1572] = 8'h33;totalMemory[1573] = 8'h2d;totalMemory[1574] = 8'h1d;totalMemory[1575] = 8'h3e;totalMemory[1576] = 8'h37;totalMemory[1577] = 8'h26;totalMemory[1578] = 8'h4b;totalMemory[1579] = 8'h41;totalMemory[1580] = 8'h30;totalMemory[1581] = 8'h62;totalMemory[1582] = 8'h56;totalMemory[1583] = 8'h46;totalMemory[1584] = 8'h7e;totalMemory[1585] = 8'h70;totalMemory[1586] = 8'h61;totalMemory[1587] = 8'h99;totalMemory[1588] = 8'h88;totalMemory[1589] = 8'h7a;totalMemory[1590] = 8'hba;totalMemory[1591] = 8'ha7;totalMemory[1592] = 8'h9a;totalMemory[1593] = 8'hd9;totalMemory[1594] = 8'hc3;totalMemory[1595] = 8'hba;totalMemory[1596] = 8'he3;totalMemory[1597] = 8'hcb;totalMemory[1598] = 8'hc4;totalMemory[1599] = 8'hea;totalMemory[1600] = 8'hd0;totalMemory[1601] = 8'hca;totalMemory[1602] = 8'hf6;totalMemory[1603] = 8'hdf;totalMemory[1604] = 8'hda;totalMemory[1605] = 8'hfb;totalMemory[1606] = 8'he5;totalMemory[1607] = 8'hdf;totalMemory[1608] = 8'he2;totalMemory[1609] = 8'hca;totalMemory[1610] = 8'hbf;totalMemory[1611] = 8'hc1;totalMemory[1612] = 8'ha6;totalMemory[1613] = 8'h94;totalMemory[1614] = 8'hc0;totalMemory[1615] = 8'ha5;totalMemory[1616] = 8'h8a;totalMemory[1617] = 8'hd2;totalMemory[1618] = 8'hb9;totalMemory[1619] = 8'h94;totalMemory[1620] = 8'hcf;totalMemory[1621] = 8'hba;totalMemory[1622] = 8'h90;totalMemory[1623] = 8'had;totalMemory[1624] = 8'h9f;totalMemory[1625] = 8'h76;totalMemory[1626] = 8'h85;totalMemory[1627] = 8'h7b;totalMemory[1628] = 8'h52;totalMemory[1629] = 8'h62;totalMemory[1630] = 8'h59;totalMemory[1631] = 8'h33;totalMemory[1632] = 8'h51;totalMemory[1633] = 8'h4a;totalMemory[1634] = 8'h21;totalMemory[1635] = 8'h51;totalMemory[1636] = 8'h4b;totalMemory[1637] = 8'h1f;totalMemory[1638] = 8'h59;totalMemory[1639] = 8'h54;totalMemory[1640] = 8'h20;totalMemory[1641] = 8'h66;totalMemory[1642] = 8'h65;totalMemory[1643] = 8'h23;totalMemory[1644] = 8'h79;totalMemory[1645] = 8'h78;totalMemory[1646] = 8'h28;totalMemory[1647] = 8'h8e;totalMemory[1648] = 8'h88;totalMemory[1649] = 8'h28;totalMemory[1650] = 8'h9f;totalMemory[1651] = 8'h93;totalMemory[1652] = 8'h25;totalMemory[1653] = 8'ha5;totalMemory[1654] = 8'h93;totalMemory[1655] = 8'h19;totalMemory[1656] = 8'ha3;totalMemory[1657] = 8'h8f;totalMemory[1658] = 8'hb;totalMemory[1659] = 8'ha6;totalMemory[1660] = 8'h90;totalMemory[1661] = 8'h6;totalMemory[1662] = 8'ha7;totalMemory[1663] = 8'h93;totalMemory[1664] = 8'hd;totalMemory[1665] = 8'h9d;totalMemory[1666] = 8'h8e;totalMemory[1667] = 8'h13;totalMemory[1668] = 8'h88;totalMemory[1669] = 8'h86;totalMemory[1670] = 8'h18;totalMemory[1671] = 8'h76;totalMemory[1672] = 8'h86;totalMemory[1673] = 8'h25;totalMemory[1674] = 8'h6b;totalMemory[1675] = 8'h86;totalMemory[1676] = 8'h2f;totalMemory[1677] = 8'h5f;totalMemory[1678] = 8'h80;totalMemory[1679] = 8'h33;totalMemory[1680] = 8'h37;totalMemory[1681] = 8'h35;totalMemory[1682] = 8'h28;totalMemory[1683] = 8'h32;totalMemory[1684] = 8'h2e;totalMemory[1685] = 8'h21;totalMemory[1686] = 8'h2e;totalMemory[1687] = 8'h29;totalMemory[1688] = 8'h1a;totalMemory[1689] = 8'h3a;totalMemory[1690] = 8'h34;totalMemory[1691] = 8'h21;totalMemory[1692] = 8'h54;totalMemory[1693] = 8'h4b;totalMemory[1694] = 8'h38;totalMemory[1695] = 8'h70;totalMemory[1696] = 8'h63;totalMemory[1697] = 8'h52;totalMemory[1698] = 8'h90;totalMemory[1699] = 8'h7f;totalMemory[1700] = 8'h70;totalMemory[1701] = 8'hb2;totalMemory[1702] = 8'h9e;totalMemory[1703] = 8'h93;totalMemory[1704] = 8'hcb;totalMemory[1705] = 8'hb6;totalMemory[1706] = 8'had;totalMemory[1707] = 8'hdd;totalMemory[1708] = 8'hc6;totalMemory[1709] = 8'hbf;totalMemory[1710] = 8'he8;totalMemory[1711] = 8'hd0;totalMemory[1712] = 8'hcb;totalMemory[1713] = 8'hf3;totalMemory[1714] = 8'hd8;totalMemory[1715] = 8'hd6;totalMemory[1716] = 8'hf6;totalMemory[1717] = 8'hdc;totalMemory[1718] = 8'hdb;totalMemory[1719] = 8'hf5;totalMemory[1720] = 8'hdb;totalMemory[1721] = 8'hd8;totalMemory[1722] = 8'hfa;totalMemory[1723] = 8'he1;totalMemory[1724] = 8'hdc;totalMemory[1725] = 8'hf9;totalMemory[1726] = 8'hdf;totalMemory[1727] = 8'hda;totalMemory[1728] = 8'he4;totalMemory[1729] = 8'hca;totalMemory[1730] = 8'hc4;totalMemory[1731] = 8'hda;totalMemory[1732] = 8'hc2;totalMemory[1733] = 8'hb9;totalMemory[1734] = 8'hdf;totalMemory[1735] = 8'hca;totalMemory[1736] = 8'hbc;totalMemory[1737] = 8'hd1;totalMemory[1738] = 8'hbf;totalMemory[1739] = 8'hab;totalMemory[1740] = 8'ha2;totalMemory[1741] = 8'h96;totalMemory[1742] = 8'h7c;totalMemory[1743] = 8'h69;totalMemory[1744] = 8'h63;totalMemory[1745] = 8'h45;totalMemory[1746] = 8'h49;totalMemory[1747] = 8'h46;totalMemory[1748] = 8'h25;totalMemory[1749] = 8'h46;totalMemory[1750] = 8'h41;totalMemory[1751] = 8'h1f;totalMemory[1752] = 8'h4c;totalMemory[1753] = 8'h47;totalMemory[1754] = 8'h21;totalMemory[1755] = 8'h58;totalMemory[1756] = 8'h52;totalMemory[1757] = 8'h24;totalMemory[1758] = 8'h6c;totalMemory[1759] = 8'h66;totalMemory[1760] = 8'h29;totalMemory[1761] = 8'h84;totalMemory[1762] = 8'h7b;totalMemory[1763] = 8'h2c;totalMemory[1764] = 8'h94;totalMemory[1765] = 8'h8b;totalMemory[1766] = 8'h2b;totalMemory[1767] = 8'h9e;totalMemory[1768] = 8'h92;totalMemory[1769] = 8'h26;totalMemory[1770] = 8'h9f;totalMemory[1771] = 8'h8f;totalMemory[1772] = 8'h1a;totalMemory[1773] = 8'h9b;totalMemory[1774] = 8'h89;totalMemory[1775] = 8'he;totalMemory[1776] = 8'h9e;totalMemory[1777] = 8'h8a;totalMemory[1778] = 8'hc;totalMemory[1779] = 8'ha4;totalMemory[1780] = 8'h90;totalMemory[1781] = 8'h11;totalMemory[1782] = 8'h9d;totalMemory[1783] = 8'h8e;totalMemory[1784] = 8'h16;totalMemory[1785] = 8'h8a;totalMemory[1786] = 8'h85;totalMemory[1787] = 8'h1b;totalMemory[1788] = 8'h76;totalMemory[1789] = 8'h7f;totalMemory[1790] = 8'h20;totalMemory[1791] = 8'h6b;totalMemory[1792] = 8'h82;totalMemory[1793] = 8'h2c;totalMemory[1794] = 8'h62;totalMemory[1795] = 8'h81;totalMemory[1796] = 8'h34;totalMemory[1797] = 8'h5a;totalMemory[1798] = 8'h7d;totalMemory[1799] = 8'h36;totalMemory[1800] = 8'h33;totalMemory[1801] = 8'h2f;totalMemory[1802] = 8'h22;totalMemory[1803] = 8'h32;totalMemory[1804] = 8'h2c;totalMemory[1805] = 8'h20;totalMemory[1806] = 8'h43;totalMemory[1807] = 8'h3b;totalMemory[1808] = 8'h2d;totalMemory[1809] = 8'h6d;totalMemory[1810] = 8'h63;totalMemory[1811] = 8'h52;totalMemory[1812] = 8'h95;totalMemory[1813] = 8'h88;totalMemory[1814] = 8'h77;totalMemory[1815] = 8'hb3;totalMemory[1816] = 8'ha0;totalMemory[1817] = 8'h93;totalMemory[1818] = 8'hd1;totalMemory[1819] = 8'hbc;totalMemory[1820] = 8'hb1;totalMemory[1821] = 8'he7;totalMemory[1822] = 8'hcf;totalMemory[1823] = 8'hc7;totalMemory[1824] = 8'hee;totalMemory[1825] = 8'hd4;totalMemory[1826] = 8'hd0;totalMemory[1827] = 8'hf3;totalMemory[1828] = 8'hd8;totalMemory[1829] = 8'hd7;totalMemory[1830] = 8'hf5;totalMemory[1831] = 8'hdb;totalMemory[1832] = 8'hdb;totalMemory[1833] = 8'hf8;totalMemory[1834] = 8'hdd;totalMemory[1835] = 8'hdd;totalMemory[1836] = 8'hfd;totalMemory[1837] = 8'he2;totalMemory[1838] = 8'he2;totalMemory[1839] = 8'hff;totalMemory[1840] = 8'he9;totalMemory[1841] = 8'he7;totalMemory[1842] = 8'hff;totalMemory[1843] = 8'hed;totalMemory[1844] = 8'hea;totalMemory[1845] = 8'hfd;totalMemory[1846] = 8'heb;totalMemory[1847] = 8'he7;totalMemory[1848] = 8'hf4;totalMemory[1849] = 8'hdf;totalMemory[1850] = 8'hdb;totalMemory[1851] = 8'hdd;totalMemory[1852] = 8'hc9;totalMemory[1853] = 8'hc4;totalMemory[1854] = 8'hb3;totalMemory[1855] = 8'ha3;totalMemory[1856] = 8'h9a;totalMemory[1857] = 8'h7f;totalMemory[1858] = 8'h74;totalMemory[1859] = 8'h66;totalMemory[1860] = 8'h53;totalMemory[1861] = 8'h4c;totalMemory[1862] = 8'h3a;totalMemory[1863] = 8'h3e;totalMemory[1864] = 8'h3c;totalMemory[1865] = 8'h22;totalMemory[1866] = 8'h40;totalMemory[1867] = 8'h3e;totalMemory[1868] = 8'h20;totalMemory[1869] = 8'h4a;totalMemory[1870] = 8'h46;totalMemory[1871] = 8'h27;totalMemory[1872] = 8'h59;totalMemory[1873] = 8'h52;totalMemory[1874] = 8'h2d;totalMemory[1875] = 8'h71;totalMemory[1876] = 8'h69;totalMemory[1877] = 8'h38;totalMemory[1878] = 8'h8a;totalMemory[1879] = 8'h81;totalMemory[1880] = 8'h40;totalMemory[1881] = 8'h9b;totalMemory[1882] = 8'h90;totalMemory[1883] = 8'h3a;totalMemory[1884] = 8'h9e;totalMemory[1885] = 8'h91;totalMemory[1886] = 8'h2d;totalMemory[1887] = 8'h98;totalMemory[1888] = 8'h89;totalMemory[1889] = 8'h1e;totalMemory[1890] = 8'h8f;totalMemory[1891] = 8'h7f;totalMemory[1892] = 8'h10;totalMemory[1893] = 8'h92;totalMemory[1894] = 8'h81;totalMemory[1895] = 8'hf;totalMemory[1896] = 8'h9d;totalMemory[1897] = 8'h8c;totalMemory[1898] = 8'h19;totalMemory[1899] = 8'h9e;totalMemory[1900] = 8'h8e;totalMemory[1901] = 8'h1e;totalMemory[1902] = 8'h8c;totalMemory[1903] = 8'h83;totalMemory[1904] = 8'h1c;totalMemory[1905] = 8'h78;totalMemory[1906] = 8'h7a;totalMemory[1907] = 8'h20;totalMemory[1908] = 8'h6b;totalMemory[1909] = 8'h79;totalMemory[1910] = 8'h28;totalMemory[1911] = 8'h65;totalMemory[1912] = 8'h7e;totalMemory[1913] = 8'h32;totalMemory[1914] = 8'h5d;totalMemory[1915] = 8'h7e;totalMemory[1916] = 8'h37;totalMemory[1917] = 8'h57;totalMemory[1918] = 8'h7c;totalMemory[1919] = 8'h3b;totalMemory[1920] = 8'h54;totalMemory[1921] = 8'h49;totalMemory[1922] = 8'h3d;totalMemory[1923] = 8'h68;totalMemory[1924] = 8'h5b;totalMemory[1925] = 8'h4f;totalMemory[1926] = 8'h85;totalMemory[1927] = 8'h77;totalMemory[1928] = 8'h6c;totalMemory[1929] = 8'hb3;totalMemory[1930] = 8'ha3;totalMemory[1931] = 8'h98;totalMemory[1932] = 8'hd2;totalMemory[1933] = 8'hbe;totalMemory[1934] = 8'hb4;totalMemory[1935] = 8'hde;totalMemory[1936] = 8'hc6;totalMemory[1937] = 8'hc0;totalMemory[1938] = 8'hed;totalMemory[1939] = 8'hd2;totalMemory[1940] = 8'hce;totalMemory[1941] = 8'hf8;totalMemory[1942] = 8'hdc;totalMemory[1943] = 8'hda;totalMemory[1944] = 8'hfa;totalMemory[1945] = 8'he1;totalMemory[1946] = 8'he0;totalMemory[1947] = 8'hfc;totalMemory[1948] = 8'he7;totalMemory[1949] = 8'he6;totalMemory[1950] = 8'hfe;totalMemory[1951] = 8'hef;totalMemory[1952] = 8'hee;totalMemory[1953] = 8'hff;totalMemory[1954] = 8'hed;totalMemory[1955] = 8'hec;totalMemory[1956] = 8'hff;totalMemory[1957] = 8'he5;totalMemory[1958] = 8'he5;totalMemory[1959] = 8'hfe;totalMemory[1960] = 8'he6;totalMemory[1961] = 8'he6;totalMemory[1962] = 8'hfc;totalMemory[1963] = 8'heb;totalMemory[1964] = 8'he8;totalMemory[1965] = 8'hf1;totalMemory[1966] = 8'he4;totalMemory[1967] = 8'hdf;totalMemory[1968] = 8'hd7;totalMemory[1969] = 8'hc8;totalMemory[1970] = 8'hc2;totalMemory[1971] = 8'ha0;totalMemory[1972] = 8'h92;totalMemory[1973] = 8'h8a;totalMemory[1974] = 8'h61;totalMemory[1975] = 8'h57;totalMemory[1976] = 8'h4d;totalMemory[1977] = 8'h3d;totalMemory[1978] = 8'h37;totalMemory[1979] = 8'h26;totalMemory[1980] = 8'h3b;totalMemory[1981] = 8'h37;totalMemory[1982] = 8'h20;totalMemory[1983] = 8'h53;totalMemory[1984] = 8'h4e;totalMemory[1985] = 8'h34;totalMemory[1986] = 8'h68;totalMemory[1987] = 8'h61;totalMemory[1988] = 8'h44;totalMemory[1989] = 8'h72;totalMemory[1990] = 8'h68;totalMemory[1991] = 8'h4b;totalMemory[1992] = 8'h85;totalMemory[1993] = 8'h79;totalMemory[1994] = 8'h54;totalMemory[1995] = 8'h9a;totalMemory[1996] = 8'h8d;totalMemory[1997] = 8'h5b;totalMemory[1998] = 8'ha1;totalMemory[1999] = 8'h94;totalMemory[2000] = 8'h52;totalMemory[2001] = 8'h9a;totalMemory[2002] = 8'h8e;totalMemory[2003] = 8'h3c;totalMemory[2004] = 8'h8e;totalMemory[2005] = 8'h83;totalMemory[2006] = 8'h28;totalMemory[2007] = 8'h82;totalMemory[2008] = 8'h79;totalMemory[2009] = 8'h1c;totalMemory[2010] = 8'h81;totalMemory[2011] = 8'h77;totalMemory[2012] = 8'h1a;totalMemory[2013] = 8'h8d;totalMemory[2014] = 8'h80;totalMemory[2015] = 8'h20;totalMemory[2016] = 8'h93;totalMemory[2017] = 8'h87;totalMemory[2018] = 8'h26;totalMemory[2019] = 8'h8c;totalMemory[2020] = 8'h83;totalMemory[2021] = 8'h27;totalMemory[2022] = 8'h79;totalMemory[2023] = 8'h78;totalMemory[2024] = 8'h22;totalMemory[2025] = 8'h6b;totalMemory[2026] = 8'h74;totalMemory[2027] = 8'h25;totalMemory[2028] = 8'h64;totalMemory[2029] = 8'h76;totalMemory[2030] = 8'h2d;totalMemory[2031] = 8'h60;totalMemory[2032] = 8'h7b;totalMemory[2033] = 8'h36;totalMemory[2034] = 8'h5c;totalMemory[2035] = 8'h7d;totalMemory[2036] = 8'h3d;totalMemory[2037] = 8'h58;totalMemory[2038] = 8'h7d;totalMemory[2039] = 8'h43;totalMemory[2040] = 8'ha7;totalMemory[2041] = 8'h97;totalMemory[2042] = 8'h8e;totalMemory[2043] = 8'hbe;totalMemory[2044] = 8'had;totalMemory[2045] = 8'ha3;totalMemory[2046] = 8'hcb;totalMemory[2047] = 8'hb8;totalMemory[2048] = 8'hb1;totalMemory[2049] = 8'hdf;totalMemory[2050] = 8'hc9;totalMemory[2051] = 8'hc4;totalMemory[2052] = 8'hef;totalMemory[2053] = 8'hd9;totalMemory[2054] = 8'hd6;totalMemory[2055] = 8'hf6;totalMemory[2056] = 8'hdf;totalMemory[2057] = 8'hde;totalMemory[2058] = 8'hf9;totalMemory[2059] = 8'hdf;totalMemory[2060] = 8'hdf;totalMemory[2061] = 8'hfb;totalMemory[2062] = 8'hdf;totalMemory[2063] = 8'hdf;totalMemory[2064] = 8'hfc;totalMemory[2065] = 8'he3;totalMemory[2066] = 8'he4;totalMemory[2067] = 8'hfd;totalMemory[2068] = 8'he8;totalMemory[2069] = 8'he9;totalMemory[2070] = 8'hfe;totalMemory[2071] = 8'hee;totalMemory[2072] = 8'hef;totalMemory[2073] = 8'hfe;totalMemory[2074] = 8'hee;totalMemory[2075] = 8'hee;totalMemory[2076] = 8'hfe;totalMemory[2077] = 8'he8;totalMemory[2078] = 8'he8;totalMemory[2079] = 8'hf5;totalMemory[2080] = 8'hdc;totalMemory[2081] = 8'hdc;totalMemory[2082] = 8'hd7;totalMemory[2083] = 8'hc0;totalMemory[2084] = 8'hbd;totalMemory[2085] = 8'haa;totalMemory[2086] = 8'h98;totalMemory[2087] = 8'h92;totalMemory[2088] = 8'h79;totalMemory[2089] = 8'h6b;totalMemory[2090] = 8'h62;totalMemory[2091] = 8'h4c;totalMemory[2092] = 8'h41;totalMemory[2093] = 8'h37;totalMemory[2094] = 8'h35;totalMemory[2095] = 8'h2c;totalMemory[2096] = 8'h1e;totalMemory[2097] = 8'h37;totalMemory[2098] = 8'h31;totalMemory[2099] = 8'h1f;totalMemory[2100] = 8'h5b;totalMemory[2101] = 8'h54;totalMemory[2102] = 8'h3f;totalMemory[2103] = 8'h96;totalMemory[2104] = 8'h8c;totalMemory[2105] = 8'h75;totalMemory[2106] = 8'hbc;totalMemory[2107] = 8'hb0;totalMemory[2108] = 8'h98;totalMemory[2109] = 8'hc1;totalMemory[2110] = 8'hb3;totalMemory[2111] = 8'h9c;totalMemory[2112] = 8'hbb;totalMemory[2113] = 8'hab;totalMemory[2114] = 8'h8f;totalMemory[2115] = 8'ha6;totalMemory[2116] = 8'h99;totalMemory[2117] = 8'h6e;totalMemory[2118] = 8'h8a;totalMemory[2119] = 8'h7f;totalMemory[2120] = 8'h46;totalMemory[2121] = 8'h77;totalMemory[2122] = 8'h6e;totalMemory[2123] = 8'h2a;totalMemory[2124] = 8'h6b;totalMemory[2125] = 8'h64;totalMemory[2126] = 8'h1a;totalMemory[2127] = 8'h6a;totalMemory[2128] = 8'h64;totalMemory[2129] = 8'h1b;totalMemory[2130] = 8'h79;totalMemory[2131] = 8'h73;totalMemory[2132] = 8'h2a;totalMemory[2133] = 8'h87;totalMemory[2134] = 8'h7e;totalMemory[2135] = 8'h33;totalMemory[2136] = 8'h86;totalMemory[2137] = 8'h7e;totalMemory[2138] = 8'h32;totalMemory[2139] = 8'h7f;totalMemory[2140] = 8'h7c;totalMemory[2141] = 8'h31;totalMemory[2142] = 8'h72;totalMemory[2143] = 8'h78;totalMemory[2144] = 8'h2e;totalMemory[2145] = 8'h68;totalMemory[2146] = 8'h76;totalMemory[2147] = 8'h30;totalMemory[2148] = 8'h60;totalMemory[2149] = 8'h77;totalMemory[2150] = 8'h33;totalMemory[2151] = 8'h5b;totalMemory[2152] = 8'h7a;totalMemory[2153] = 8'h39;totalMemory[2154] = 8'h5a;totalMemory[2155] = 8'h7d;totalMemory[2156] = 8'h40;totalMemory[2157] = 8'h5a;totalMemory[2158] = 8'h7f;totalMemory[2159] = 8'h49;totalMemory[2160] = 8'he0;totalMemory[2161] = 8'hcb;totalMemory[2162] = 8'hc9;totalMemory[2163] = 8'hea;totalMemory[2164] = 8'hd5;totalMemory[2165] = 8'hd4;totalMemory[2166] = 8'hec;totalMemory[2167] = 8'hd6;totalMemory[2168] = 8'hd5;totalMemory[2169] = 8'hf2;totalMemory[2170] = 8'hdb;totalMemory[2171] = 8'hdb;totalMemory[2172] = 8'hfa;totalMemory[2173] = 8'he5;totalMemory[2174] = 8'he6;totalMemory[2175] = 8'hfe;totalMemory[2176] = 8'hea;totalMemory[2177] = 8'hec;totalMemory[2178] = 8'hfd;totalMemory[2179] = 8'he6;totalMemory[2180] = 8'he8;totalMemory[2181] = 8'hfb;totalMemory[2182] = 8'he1;totalMemory[2183] = 8'he4;totalMemory[2184] = 8'hfb;totalMemory[2185] = 8'he1;totalMemory[2186] = 8'he4;totalMemory[2187] = 8'hfa;totalMemory[2188] = 8'he0;totalMemory[2189] = 8'he2;totalMemory[2190] = 8'hf8;totalMemory[2191] = 8'he0;totalMemory[2192] = 8'he2;totalMemory[2193] = 8'hf7;totalMemory[2194] = 8'he0;totalMemory[2195] = 8'he3;totalMemory[2196] = 8'hec;totalMemory[2197] = 8'hd7;totalMemory[2198] = 8'hd9;totalMemory[2199] = 8'hc4;totalMemory[2200] = 8'hb0;totalMemory[2201] = 8'haf;totalMemory[2202] = 8'h84;totalMemory[2203] = 8'h73;totalMemory[2204] = 8'h6e;totalMemory[2205] = 8'h4f;totalMemory[2206] = 8'h42;totalMemory[2207] = 8'h38;totalMemory[2208] = 8'h35;totalMemory[2209] = 8'h2a;totalMemory[2210] = 8'h1e;totalMemory[2211] = 8'h31;totalMemory[2212] = 8'h26;totalMemory[2213] = 8'h17;totalMemory[2214] = 8'h42;totalMemory[2215] = 8'h36;totalMemory[2216] = 8'h25;totalMemory[2217] = 8'h68;totalMemory[2218] = 8'h5b;totalMemory[2219] = 8'h49;totalMemory[2220] = 8'h96;totalMemory[2221] = 8'h87;totalMemory[2222] = 8'h77;totalMemory[2223] = 8'hc3;totalMemory[2224] = 8'hb2;totalMemory[2225] = 8'ha4;totalMemory[2226] = 8'he6;totalMemory[2227] = 8'hd5;totalMemory[2228] = 8'hc8;totalMemory[2229] = 8'hec;totalMemory[2230] = 8'hdc;totalMemory[2231] = 8'hd0;totalMemory[2232] = 8'hc0;totalMemory[2233] = 8'hb4;totalMemory[2234] = 8'ha4;totalMemory[2235] = 8'h7d;totalMemory[2236] = 8'h75;totalMemory[2237] = 8'h5c;totalMemory[2238] = 8'h52;totalMemory[2239] = 8'h4d;totalMemory[2240] = 8'h2b;totalMemory[2241] = 8'h46;totalMemory[2242] = 8'h43;totalMemory[2243] = 8'h18;totalMemory[2244] = 8'h4e;totalMemory[2245] = 8'h4a;totalMemory[2246] = 8'h1b;totalMemory[2247] = 8'h6a;totalMemory[2248] = 8'h64;totalMemory[2249] = 8'h34;totalMemory[2250] = 8'h86;totalMemory[2251] = 8'h80;totalMemory[2252] = 8'h4e;totalMemory[2253] = 8'h8f;totalMemory[2254] = 8'h89;totalMemory[2255] = 8'h54;totalMemory[2256] = 8'h86;totalMemory[2257] = 8'h82;totalMemory[2258] = 8'h4a;totalMemory[2259] = 8'h7a;totalMemory[2260] = 8'h7c;totalMemory[2261] = 8'h3d;totalMemory[2262] = 8'h6f;totalMemory[2263] = 8'h7a;totalMemory[2264] = 8'h36;totalMemory[2265] = 8'h67;totalMemory[2266] = 8'h7a;totalMemory[2267] = 8'h36;totalMemory[2268] = 8'h62;totalMemory[2269] = 8'h7c;totalMemory[2270] = 8'h3a;totalMemory[2271] = 8'h5c;totalMemory[2272] = 8'h7e;totalMemory[2273] = 8'h3e;totalMemory[2274] = 8'h57;totalMemory[2275] = 8'h7e;totalMemory[2276] = 8'h42;totalMemory[2277] = 8'h57;totalMemory[2278] = 8'h7f;totalMemory[2279] = 8'h4a;totalMemory[2280] = 8'hef;totalMemory[2281] = 8'hd9;totalMemory[2282] = 8'hdb;totalMemory[2283] = 8'hf4;totalMemory[2284] = 8'hdd;totalMemory[2285] = 8'he0;totalMemory[2286] = 8'hf7;totalMemory[2287] = 8'hdf;totalMemory[2288] = 8'he2;totalMemory[2289] = 8'hf9;totalMemory[2290] = 8'he1;totalMemory[2291] = 8'he4;totalMemory[2292] = 8'hfa;totalMemory[2293] = 8'he3;totalMemory[2294] = 8'he6;totalMemory[2295] = 8'hf9;totalMemory[2296] = 8'he4;totalMemory[2297] = 8'he7;totalMemory[2298] = 8'hf9;totalMemory[2299] = 8'he4;totalMemory[2300] = 8'he6;totalMemory[2301] = 8'hfa;totalMemory[2302] = 8'he5;totalMemory[2303] = 8'he7;totalMemory[2304] = 8'hf8;totalMemory[2305] = 8'he1;totalMemory[2306] = 8'he3;totalMemory[2307] = 8'hf2;totalMemory[2308] = 8'hdc;totalMemory[2309] = 8'hde;totalMemory[2310] = 8'hea;totalMemory[2311] = 8'hd6;totalMemory[2312] = 8'hd7;totalMemory[2313] = 8'hd8;totalMemory[2314] = 8'hc6;totalMemory[2315] = 8'hc7;totalMemory[2316] = 8'hb1;totalMemory[2317] = 8'ha1;totalMemory[2318] = 8'ha0;totalMemory[2319] = 8'h74;totalMemory[2320] = 8'h66;totalMemory[2321] = 8'h61;totalMemory[2322] = 8'h44;totalMemory[2323] = 8'h37;totalMemory[2324] = 8'h2d;totalMemory[2325] = 8'h33;totalMemory[2326] = 8'h28;totalMemory[2327] = 8'h1b;totalMemory[2328] = 8'h40;totalMemory[2329] = 8'h35;totalMemory[2330] = 8'h24;totalMemory[2331] = 8'h5e;totalMemory[2332] = 8'h51;totalMemory[2333] = 8'h40;totalMemory[2334] = 8'h87;totalMemory[2335] = 8'h78;totalMemory[2336] = 8'h68;totalMemory[2337] = 8'hb8;totalMemory[2338] = 8'ha7;totalMemory[2339] = 8'h99;totalMemory[2340] = 8'hd2;totalMemory[2341] = 8'hbe;totalMemory[2342] = 8'hb3;totalMemory[2343] = 8'hd4;totalMemory[2344] = 8'hbf;totalMemory[2345] = 8'hb8;totalMemory[2346] = 8'hd9;totalMemory[2347] = 8'hc5;totalMemory[2348] = 8'hc0;totalMemory[2349] = 8'hca;totalMemory[2350] = 8'hb9;totalMemory[2351] = 8'hb4;totalMemory[2352] = 8'h8d;totalMemory[2353] = 8'h81;totalMemory[2354] = 8'h79;totalMemory[2355] = 8'h4f;totalMemory[2356] = 8'h49;totalMemory[2357] = 8'h3b;totalMemory[2358] = 8'h37;totalMemory[2359] = 8'h34;totalMemory[2360] = 8'h1f;totalMemory[2361] = 8'h36;totalMemory[2362] = 8'h34;totalMemory[2363] = 8'h1a;totalMemory[2364] = 8'h59;totalMemory[2365] = 8'h56;totalMemory[2366] = 8'h39;totalMemory[2367] = 8'h8c;totalMemory[2368] = 8'h86;totalMemory[2369] = 8'h68;totalMemory[2370] = 8'ha2;totalMemory[2371] = 8'h9b;totalMemory[2372] = 8'h7c;totalMemory[2373] = 8'ha1;totalMemory[2374] = 8'h9b;totalMemory[2375] = 8'h7a;totalMemory[2376] = 8'h8e;totalMemory[2377] = 8'h8d;totalMemory[2378] = 8'h64;totalMemory[2379] = 8'h78;totalMemory[2380] = 8'h7f;totalMemory[2381] = 8'h48;totalMemory[2382] = 8'h6a;totalMemory[2383] = 8'h7a;totalMemory[2384] = 8'h3b;totalMemory[2385] = 8'h63;totalMemory[2386] = 8'h7a;totalMemory[2387] = 8'h39;totalMemory[2388] = 8'h5d;totalMemory[2389] = 8'h7b;totalMemory[2390] = 8'h3a;totalMemory[2391] = 8'h59;totalMemory[2392] = 8'h7e;totalMemory[2393] = 8'h3d;totalMemory[2394] = 8'h57;totalMemory[2395] = 8'h80;totalMemory[2396] = 8'h44;totalMemory[2397] = 8'h58;totalMemory[2398] = 8'h82;totalMemory[2399] = 8'h4a;
end
  
  always @(start) begin
    if (start == 1'b1) begin
      // Read image hex value into temporary varibale
      for (i = 0; i < WIDTH * HEIGHT * 3; i = i + 1) begin
        tempBMP[i] = totalMemory[i][7:0];
      end

      // Matlab script to convert from bitmap image to hex process from the last row to the first row, so the verilog code need to operate the same.
      for (i = 0; i < HEIGHT; i = i + 1) begin
        for (j = 0; j < WIDTH; j = j + 1) begin
          tempRedValue[WIDTH*i+j]   = tempBMP[WIDTH*3*(HEIGHT-i-1)+3*j+0];
          tempGreenValue[WIDTH*i+j] = tempBMP[WIDTH*3*(HEIGHT-i-1)+3*j+1];
          tempBlueValue[WIDTH*i+j]  = tempBMP[WIDTH*3*(HEIGHT-i-1)+3*j+2];
        end
      end
    end
  end

  //--- BEGIN TO READ IMAGE FILE ONCE RESET WAS HIGH ---

  always @(posedge HCLK, negedge HRESET) begin
    if (!HRESET) begin
      start <= 0;
      HRESETDelay <= 0;
    end else begin
      HRESETDelay <= HRESET;
      if (HRESET == 1'b1 && HRESETDelay == 1'b0) start <= 1'b1;
      //else start <= 1'b0;
    end
  end

  /*--- FSM for reading RGB888 data from memory ---
    --- Creating hsync and vsync pulse --- */

  always @(posedge HCLK, negedge HRESET) begin
    if (~HRESET) currentState <= ST_IDLE;
    else currentState <= nextState;
  end

  //--- State transition ---

  always @(*) begin
    case (currentState)
      ST_IDLE: begin
        if (start) nextState = ST_VSYNC;
        else nextState = ST_IDLE;
      end
      ST_VSYNC: begin
        if (vsyncControlCounter == STARTUP_DELAY) nextState = ST_HSYNC;
        else nextState = ST_VSYNC;
      end
      ST_HSYNC: begin
        if (hsyncControlCounter == HSYNC_DELAY) nextState = ST_DATA;
        else nextState = ST_HSYNC;
      end
      ST_DATA: begin
        if (ctrl_done) nextState = ST_IDLE;
        else begin
          if (colIndex == WIDTH - 2) nextState = ST_HSYNC;
          else nextState = ST_DATA;
        end
      end
    endcase
  end

  //--- Counting for time period of vsync, hsync, data processing ---

  always @(*) begin
    vsyncControlSignal = 0;
    hsyncControlSignal = 0;
    dataProcessingControlSignal = 0;

    case (currentState)
      ST_VSYNC: vsyncControlSignal = 1;
      ST_HSYNC: hsyncControlSignal = 1;
      ST_DATA:  dataProcessingControlSignal = 1;
    endcase
  end

  // Counter for vsync, hsync
  always @(posedge HCLK, negedge HRESET) begin
    begin
      if (~HRESET) begin
        vsyncControlCounter <= 0;
        hsyncControlCounter <= 0;
      end else begin
        if (vsyncControlSignal) vsyncControlCounter <= vsyncControlCounter + 1;
        else vsyncControlCounter <= 0;
        if (hsyncControlSignal) hsyncControlCounter <= hsyncControlCounter + 1;
        else hsyncControlCounter <= 0;
      end
    end
  end

  // Counting column and row index for reading memory
  always @(posedge HCLK, negedge HRESET) begin
    if (~HRESET) begin
      rowIndex <= 0;
      colIndex <= 0;
    end else begin
      if (dataProcessingControlSignal) begin
        if (colIndex == WIDTH - 2) begin
          rowIndex <= rowIndex + 1;
          colIndex <= 0;
        end else colIndex <= colIndex + 2;  // Reading 2 pixels in parallel
      end
    end
  end

  //--- Data counting ---

  always @(posedge HCLK, negedge HRESET) begin
    if (~HRESET) pixelDataCount <= 0;
    else begin
      if (dataProcessingControlSignal) pixelDataCount <= pixelDataCount + 1;
    end
  end

  assign VSYNC = vsyncControlSignal;
  assign ctrl_done = (pixelDataCount == WIDTH * HEIGHT / 2 - 1) ? 1'b1 : 1'b0;

  //--- Image processing ---

  always @(posedge HCLK) begin
    HSYNC   = 1'b0;
    DATA_R0 = 0;
    DATA_G0 = 0;
    DATA_B0 = 0;
    DATA_R1 = 0;
    DATA_G1 = 0;
    DATA_B1 = 0;

    if (dataProcessingControlSignal) begin
      HSYNC = 1'b1;
      // BRIGHTNESS ADDING OPERATION
      if (increaseBrightness == 1'b1) begin
        tempConBriR0 = tempRedValue[WIDTH*rowIndex+colIndex] + BRIGHTNESS_VALUE;
        if (tempConBriR0 > 255) DATA_R0 = 255;
        else DATA_R0 = tempRedValue[WIDTH*rowIndex+colIndex] + BRIGHTNESS_VALUE;

        tempConBriR1 = tempRedValue[WIDTH*rowIndex+colIndex+1] + BRIGHTNESS_VALUE;
        if (tempConBriR1 > 255) DATA_R1 = 255;
        else DATA_R1 = tempRedValue[WIDTH*rowIndex+colIndex+1] + BRIGHTNESS_VALUE;

        tempConBriG0 = tempGreenValue[WIDTH*rowIndex+colIndex] + BRIGHTNESS_VALUE;
        if (tempConBriG0 > 255) DATA_G0 = 255;
        else DATA_G0 = tempGreenValue[WIDTH*rowIndex+colIndex] + BRIGHTNESS_VALUE;

        tempConBriG1 = tempGreenValue[WIDTH*rowIndex+colIndex+1] + BRIGHTNESS_VALUE;
        if (tempConBriG1 > 255) DATA_G1 = 255;
        else DATA_G1 = tempGreenValue[WIDTH*rowIndex+colIndex+1] + BRIGHTNESS_VALUE;

        tempConBriB0 = tempBlueValue[WIDTH*rowIndex+colIndex] + BRIGHTNESS_VALUE;
        if (tempConBriB0 > 255) DATA_B0 = 255;
        else DATA_B0 = tempBlueValue[WIDTH*rowIndex+colIndex] + BRIGHTNESS_VALUE;

        tempConBriB1 = tempBlueValue[WIDTH*rowIndex+colIndex+1] + BRIGHTNESS_VALUE;
        if (tempConBriB1 > 255) DATA_B1 = 255;
        else DATA_B1 = tempBlueValue[WIDTH*rowIndex+colIndex+1] + BRIGHTNESS_VALUE;
      end  // BRIGHTNESS SUBTRACTION OPERATION
      else if (decreaseBrightness == 1'b1) begin
        tempConBriR0 = tempRedValue[WIDTH*rowIndex+colIndex] - BRIGHTNESS_VALUE;
        if (tempConBriR0 < 0) DATA_R0 = 0;
        else DATA_R0 = tempRedValue[WIDTH*rowIndex+colIndex] - BRIGHTNESS_VALUE;

        tempConBriR1 = tempRedValue[WIDTH*rowIndex+colIndex+1] - BRIGHTNESS_VALUE;
        if (tempConBriR1 < 0) DATA_R1 = 0;
        else DATA_R1 = tempRedValue[WIDTH*rowIndex+colIndex+1] - BRIGHTNESS_VALUE;

        tempConBriG0 = tempGreenValue[WIDTH*rowIndex+colIndex] - BRIGHTNESS_VALUE;
        if (tempConBriG0 < 0) DATA_G0 = 0;
        else DATA_G0 = tempGreenValue[WIDTH*rowIndex+colIndex] - BRIGHTNESS_VALUE;

        tempConBriG1 = tempGreenValue[WIDTH*rowIndex+colIndex+1] - BRIGHTNESS_VALUE;
        if (tempConBriG1 < 0) DATA_G1 = 0;
        else DATA_G1 = tempGreenValue[WIDTH*rowIndex+colIndex+1] - BRIGHTNESS_VALUE;

        tempConBriB0 = tempBlueValue[WIDTH*rowIndex+colIndex] - BRIGHTNESS_VALUE;
        if (tempConBriB0 < 0) DATA_B0 = 0;
        else DATA_B0 = tempBlueValue[WIDTH*rowIndex+colIndex] - BRIGHTNESS_VALUE;

        tempConBriB1 = tempBlueValue[WIDTH*rowIndex+colIndex+1] - BRIGHTNESS_VALUE;
        if (tempConBriB1 < 0) DATA_B1 = 0;
        else DATA_B1 = tempBlueValue[WIDTH*rowIndex+colIndex+1] - BRIGHTNESS_VALUE;
      end else if (invert == 1'b1) begin
        tempInvThre2 = (tempRedValue[WIDTH*rowIndex+colIndex] + tempGreenValue[WIDTH*rowIndex+colIndex] + tempBlueValue[WIDTH*rowIndex+colIndex]) / 3;
        DATA_R0 = 255 - tempInvThre2;
        DATA_G0 = 255 - tempInvThre2;
        DATA_B0 = 255 - tempInvThre2;

        tempInvThre4 = (tempRedValue[WIDTH*rowIndex+colIndex + 1] + tempGreenValue[WIDTH*rowIndex+colIndex + 1] + tempBlueValue[WIDTH*rowIndex+colIndex + 1]) / 3;
        DATA_R1 = 255 - tempInvThre4;
        DATA_G1 = 255 - tempInvThre4;
        DATA_B1 = 255 - tempInvThre4;
      end else if (threshold == 1'b1) begin
        tempInvThre = (tempRedValue[WIDTH*rowIndex+colIndex] + tempGreenValue[WIDTH*rowIndex+colIndex] + tempBlueValue[WIDTH*rowIndex+colIndex]) / 3;
        if (tempInvThre > THRESHOLD) begin
          DATA_R0 = 255;
          DATA_G0 = 255;
          DATA_B0 = 255;
        end else begin
          DATA_R0 = 0;
          DATA_G0 = 0;
          DATA_B0 = 0;
        end

        tempInvThre1 = (tempRedValue[WIDTH*rowIndex+colIndex+1] + tempGreenValue[WIDTH*rowIndex+colIndex+1] + tempBlueValue[WIDTH*rowIndex+colIndex+1]) / 3;
        if (tempInvThre1 > THRESHOLD) begin
          DATA_R1 = 255;
          DATA_G1 = 255;
          DATA_B1 = 255;
        end else begin
          DATA_R1 = 0;
          DATA_G1 = 0;
          DATA_B1 = 0;
        end
      end else begin
        DATA_R0 = tempRedValue[WIDTH*rowIndex+colIndex];
        DATA_R1 = tempRedValue[WIDTH*rowIndex+colIndex+1];
        DATA_G0 = tempGreenValue[WIDTH*rowIndex+colIndex];
        DATA_G1 = tempGreenValue[WIDTH*rowIndex+colIndex+1];
        DATA_B0 = tempBlueValue[WIDTH*rowIndex+colIndex];
        DATA_B1 = tempBlueValue[WIDTH*rowIndex+colIndex+1];
      end
    end
  end

endmodule
