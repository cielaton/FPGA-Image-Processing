module FPGA_Image_Processing (input clk);
endmodule